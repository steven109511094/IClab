`ifdef RTL
    `define CYCLE_TIME 20
    `define RTL_GATE
`elsif GATE
    `define CYCLE_TIME 20
    `define RTL_GATE
`elsif CHIP
    `define CYCLE_TIME 20
    `define CHIP_POST 
`elsif POST
    `define CYCLE_TIME 20
    `define CHIP_POST 
`endif


`ifdef FUNC
`define MAX_WAIT_READY_CYCLE 2000
`endif
`ifdef PERF
`define MAX_WAIT_READY_CYCLE 100000
`endif


`include "../00_TESTBED/MEM_MAP_define.v"
`include "../00_TESTBED/pseudo_DRAM_data.v"
`include "../00_TESTBED/pseudo_DRAM_inst.v"

module PATTERN
`protected
3(,+(5]N_TbUJ+0K<#URQW&].5Wc,-5E/;BZ?E#cM4gHD+,QJ0-b+)JCS4B05]02
d()]ODf98I1N(KBEN+LE&_WP>e(B@/3PLM((E:209#UTWAO-W7XN260+S0U#XMgN
;DKYF9S03](#8WKNZ7Q48(K7,b<2V/R_V)W2WbD\4CT?WS&3UPJWE\PWf-g=c2dJ
.&ecO6?.@CR<<ZV/CSP.\^/@Ld&0@K5+9379,XWT5RS4?_M,FU?4T-@N+HL?e<Yb
@gN0aJLY^\_:/Wg&XZa]9(&-24G?6R>g+fJIM2BPB+,AA3NgA^+.P,d7DJYfPLO,
A3:[Z+R+;?BPWP=)V)(7LW:3P[B_@C804J&E:_[g22ZYfUMX?23E]a+H&]:X@HGP
IIIQ8>DP.[2K_5:6NHXG,WST_;,1b>2=M(ZER/4UP)>UdSA9,>C4TLd+8/N)/#B6
H9T=0VDN/c,&0;VeH[TAHa2a4?H9b[M3T(3=3+]SL[UZE#2#^GgcBB50J<R&CX=F
[+R]LXbC,:/eGOR(7M8b0_K)3(<//SPVYTf6KbE&12^-&6_8[g<PH,D.aP93aJ<g
N7SS^W0MSY@@WOFOM9/a8SFI>g>X?3eKf-?d<8_/NS-@/Oc:g:4GTTD2F;_PUJKH
6?98d(,dBTf3g5c)81@4JT9?f<N(F<[-Rb?-CORUN6C>62#BO&e8?BFa8;=aacOf
?L?UG&fVD2PTd6A>PZGD1^7#3^fcWgg._bCG)@HDPU0<,<A@gJ</BVb]A_2Se:>f
Qg\,&-[[T=WA<L;(8VMQ[c(SNB=^JVcS;:b[P4E138Z_Q?B0+PNJ2Hfd,e>T54I?
8[.89,+NfTQaIX=07E<MKf1??9d#9?A+?#;5?)Vd238M;?MA@g8L+,:,JJZ)T3KH
6=[N@4^4T#eH2#5:/>;U6PXSW,V8f/9806\J07gM<f^I=6X(^gX\:W2dCG1#]Bbf
<AKZ_1N24H6QNGV<XV<7,H<UHC0S8J;KE[5YHa374?daN;UgG83[?6a_38)YOL@D
S/0a(PZSU(H0dJd<M6E5eKeZ\GQPA4-#0N.+?.YO=P^SYba(^cGJcD/8?Tf=N;[[
H>^/4Xg2AI5Gdb];Y,N4:Z1bYU94^J3=C[FWQJTA4+&YX@>:7O,:Pf@gAgY[XPZa
;?A\.E@5He^XD:BAK0YFTNDDYe]=5++,-P\@W3efJDI2Q[+a?9bX7DfN#/GCP/T1
X^0X<.)KM\];>-P&]GJR0&a;3YQ;=]K&6&-,6feN&;(NE,I,3W=<aBK.>RT;FW.f
-bgd,Ab38O6LgWK@]J&c^^:1_,f\09/ORMK?ZPBZ(F].GPZcA5MXJ:H9]BIS;9PR
YBMT5gTE?51b+FbMNA#CYV]^;:DOR7J)>W5)A\I:#WPcZ:6H8aW&a2gGTF9bK3:P
TH<RE=78<)eNM6.\R+OWQBYA12bdR2I@^1Ng^dd8SXRSR>?NQa;7\M5Q2f</=5XU
U1bK)c,YIHF;QJUXf[^:E5=(S<WgE^EK/cSP;_UU8+6<@T:V5>Q@G8ZWF6(N1>A@
8>>OATL@SSPFLBZEE5=RH+Y5)Ef/C(:\637H:+a535O4Y&FI_-6S#WK,<0]&<d[J
GeUfLBc.7[&:/LODW@H>3/4AcB,GfZFTTS;IQRPRL8VDf[A5JcYf;8\3/Y,9Y./f
HWQ,LVfNUHGf69_PTb@P]C+&SD+/(SPeLa+FZD)C_][\].8Hc/(Z.8>>8F_Z[YbD
b7=cDMgVR7TgK?6K_;O9QP^+OOI4T_WDC@6_c5]>#eZ1R-E\IYg>S?U<8Z4.W5SD
UJ,52e1Ua?5(J(-=b(4g&aObO=K<bQZPP-N?OS&1R1;KHEY+-,-^98ac/FF2N(I.
7A>5_5ZKLD-DI4\-L:B?Z3IedIL>:WQW:7JL8CG,&H439J?_@IW=]YTK[bT:W8I@
[2GUW5ZDPR;IJ<HIP;7[;JC?O=gFG+;FP[+7ZG\[+&(PG/Q9>VFgVf;g>.AALG:#
50ZUVIC<UUAAK#TEa9c3Y[PVUgRA&7L#92;7&eBafc\7aP\=A;X1&]aeRKQD.I/C
aAJg2QHR]C6V2XS/;-,;(AHLDPK1R>+2fQKY..\ZW8H>5.Ie9P.]]W:J3BTdXPdc
I#geNE:E3AGD[TLaZ??>WHbM@3SCI8N55]A),/JP42(W.SAE+_TM-K@I,d][#&F+
Q/f6FX/5[LK2/DY/F-LcdX\AYbY0fO+OK+X6CX-VS0Lc^B4eJ@:a#)@08T\2@_J_
)g[P/1MF.G3GdES6;CH<cRLFTa=D.1/a==2:W#2?8GF.C0G5G0gQCS8dY29Q0U/9
WBbccW.)CFL<AS5QQK@>G7=7_X\(LeFIUPULQF-/]7WO9aNZ>,P:K^JWTMECYO9>
=Z6.LbY4#N?P5fF1O2PNYD7PO.QU.>0WHW\4KZI\Ma=,.,TKAU>dB#PB5.X,-G,;
?P<>(W2\:cDNCd,3N3O5MZ>S0[^Z;P76@LMGT_WYRLHYC)N#fARcEMdRGdXXc=_-
f/^/9\WJb])LB@Y3.gfPP_JW9R(I:gAZ=61cO11DfP\Sbf:c]K6@-@e6TB/PLX+]
FVBTP8I9H@Pf-SX?Ue-+b)MJVE<^H:;IEI9S[d8^SOOd]&O47W;KWA+c^K76IL9Q
1\^dEQ2,]<,dBVFg8\41OLXR0XT^I&geTSXf3EC79-1_3:fcG+@IaCCAbH/:>/VI
O_3&@;5M#bXMW87P;)4-#ND?O:;>KaL.)P;=4@:URG&QCG3IIRS6D.X,O&MVX__d
Q2f_RJd-JV5d0.N3D(9KU]^f8A;G#TU__:IT(g]N)(67ZY(;Oca#6DQ.Pc5CP6eR
N15PU6(VGJL)&ZbP2#>^9[VX_D^+]fP&C3#X\P08A\d=&&b]46ALDZYe&2B5E(=]
<-G<gBO7Q9c-BeM)/g,b2+?dPH/H,#XaI4SP0)NY+U1]B:7a^\<58OW48^H.fR:R
HC2-56gNcE4<Zc[L4SBYBZ]\e.=E-KaG^E2:UXBP1?.-d)S9JCB<_.7WJJNY=@Zb
]d)CU@2b3Q:\EN\Xa@]W<c<M0dRf6=C5+O=\\H2R[eN,(87401&(,5M015)PCGD4
A)U+WUS[B?[YI_N(^bKgG0UJWVBW39>&b<IEe-0]/_a\:1>?aNKeEc.P:3=e-.H9
=ZdJY@J;^g2Pc@M7b_?5XB<GLb1R/G,[CO##\=Z:,17O8#U,(>2GGMYKY/_\2^BC
d>Q765c3A;+CeD_+17PVU@:8HF#cL7Y@I/2:@MA13Z1HIU[Sd=II[J5J].LFBYe:
@QO>:V,?[2S>f1&LH)M.G-MPO#;QQf1Q9>8gD.Q[g+[6c)WVONf-^I?#OBdKe5e3
e,T]MF_Kg<VgRIRHVKRcJ^,:P<bYCR\NRM?4K;]3?;.ILg75TT^?\_Y(V2R=KH9(
a+>&;X;YLdcT]W=NF09-XEL-7ND]^\b]c:33a@PK48BVg_BH[7LCA.^T-6>KHegF
PC,W-D+De9^#U48bQ2e02\eW1JO/e(Nc;4V=13>1d#X]&)aHeaBJa-&J\Q>#HSSa
6LaUJE2I/TL\:HD6V]<a<g(#B<K0XA@..fa]]C9[b\2XW^TH7X;=75@9E)<W:d7a
(RB=B(C9F]FSA@[IEP8H<6.,T#R7a?<M&Tfe;XOUca;U[cc?^Xa[8Nb#bH<;,ET#
UQOJ#?I5&K1CZdJ>M-?M]feRB4P[Le+D6(SG58?(6TWZXIfGU;8GbS9R@(M3UMF?
Y;?H4O6V,cQ)d6bC5Zfd3M@+F<4H#FbLHTebIbY?CA=W/.H-TgW7NAPJ]g\[?+]E
(c-<EDdTfN2a&P1G86_SJPH0RdMcGZ]ZY2+2AQK7&G&1aCD(/N=X)6SU,X8O^?)K
H6^4/);9Fg3a1D3UG(>23ba8CcbKTT;GaU6&/SO<\BM9D:?0b;I1AA;]2H&=f#(5
S:?L@geN^P>:5H\2JOdH87D()AUG0T3->d6L0#^>[H@FTc_\V5V_O+(ac=^cK\]9
P1H3Ld+S8Sa8&F0E,0;476:)4G9d48(6?G\_)74/>a<d@9:@\U&QH?bVXID)@E19
5-4C?#&DbLd^#A1V9D.R+W)7.gb2D<I02E>J8+SQ9>51bO]A>?\==D;51V>FM^(B
9=K@[Sg(cGOc,Q#Ob]4/#NQU/F<#KU97M8fD.QbWd:f4K(.+SSfUc(<0K=4GER0U
MCSHQ?Kf?M>R-KF_eWWX=/&M;W4<#DBD,FLOZ44XO]GT9(-AXA;WaYEa[d6c[9<S
ga^CYVJef>T,^W_;O.IN-.4G-.Q35.P9Y@Zf7V46R1ASX#V4VZI???FLILGR#d/E
,JHEGG=1;Tc<5FegQ]]L?e/0O^LS(G.CI5D98[1(?0G[M#(Y]V6WP):1)_Y\/QL9
PDXQF][GXUE5gBKK5]Q:M8dCf:]JYX3Q^^=2TKeE:&HE0C2^=)=X&?H(\-:3JYgR
8MdZH9TbCFSVIE?)U^\SM_V\7;_U2Tf;UP19)2G0)(KV39KdY>Yc(/73F/RgK6(_
E7:+KF#V[P4HO7B=[(W>TCPHNEP:GP-I&C5X7J\1BdQ&UTa^WTW:,@66Pc>S3+J4
aZ#d4,>L\W(c<28929K24WSa.DO?>ULM5<M6(9#c)LMSL3X?dKT6-8;DYbBRE_4H
1(32D.[XKD62^.U_&0JfGfZeZB@e07#gSD-C>]T/?a_D[7G:(OQ3F9gV9/0dDKQ7
XcM7g.C1a+_D\[.8YVF90TRG7I&=^S24(P#X^bC]K&f-F8:#KMNK3T)E;b67bD]?
W1Pc</DE(0-(RU.,S@N=[A7UgO@PJ[W5-NgfG)1AG-d4S#44:c[[=LeIL-,\G?N5
)/A5XSNV/>>e(P:(10_CHS+VZ(f1DeYM-J\018(I.V&,5cF84b.C[\_QI+R.dLf_
=f?M&D+.4PW)8V#Z/@2a\MdP1cB6WT9R403MGcSf(7[2D(BCe[,R=d_[L?55[eb3
YeOJ#AF.aQP#3g]c.K30A9FEWOQ>(\g.cYf_W6EY.NOaN@eeK3]14ddGJA0H:5S7
1#8D]Od5,KfQ9WM(1JU)6H-]XH(MKJ4V+Q38F^7dH,GAKc<SQ:dL)[Q+0WX<2Z((
gE4,+R76_4&J5f/VgJgEEIML4/ePG1I-0#&Bf(6@VbN7YZ?D[C\Z/[.J]6gB8HR^
?4TNe7&U42MD65]T]QPCa)UE7HF/UZCZW#7++.,c,fV;G^eFXafV]DVf_5YKH[R?
Jg/X&G>-H_#?8B\#SISSZXfcBI@&G;PaY^Q@(Y^/B[FS>@,HEA.f8LC=O@)/\1d+
/8eE&HbOR5F1#O7(?[9;5g6NY9O/#e0Q]W7=Cg@J5?V,KK7BFBJ_/1292e8)#7VW
=M?^<H67gM\>E1HdHXO;]]:7K>Y0(266eVcQR>(4L5.\@9bAPF:&992=/WP?/F9/
O:&fd\0;B@;I3-_V)0I::::d/I?R[EKd?ZUXS-X/.cTW4O,-WQ-TbE=2+\#aW?YZ
2J3(F2gJ(2PKFM8>;=>^Nd8(M_UU9Zd5GY]0#\4][]Gfcc(S@-3,>\R54QU8JF4M
SP[JOCK.2f=6+D5_cfN5VD]b5?F\/F_E_1SS,IMeWRK]&TZe)A,c]7R;QX5Z]#P0
\\8@c.)GMC+L)5J=KTU:cCg:FBQQDQBPH&V?/B\057<G:21g^5M>+/c>(1K.-38F
]#]P20AR>,WeL;.X=a^R2Q5GW6.KggW-H(#YG&Y?cBONIcdUDOe6?0\/Z;^Ue@_S
e1?BIRFCCMORZKFVba?H(I]=f?6g/?\#cd0b44@FBbMT-2P:Zg9J;,+S?#J.0F(f
9?b8\R=OD1:8UX2Qd]V<6HJ<97G,FNSNG.FGS3a71US)+8=Qa)T(OM[G],?acf7L
0YHgdD7f.aJX:+#VFJ=?<_8H^)ILJ1d/K-c>V8cNBX5F);OX]LW1=e&(I(MJ2WBb
bA#(=Db&:[I<C58IRM:K\1Y&^d<aDE(^J/?(=_UG>a]PM>^>[:/4fbP]XN)ZB>2@
P0bCdYHJC3/e--42PY^QNA>]QL:HeL0-f6:0VgX?RNLa\H]9_O7?dS+NCWdP1?eJ
C-H)cOGCWgF,OfDP46#/+5?\BKD/G<DI&Z>Mfa\(6+LA@.KV8?J=^67fcX<4YX32
^16JCO36K.^P#=+bS1f7Y+^0Ucc]2UEe5S<7,fIA;.V61L7BJf6?1;)ZF(f,Q>fW
;KGCQ(6W[fcTa3--.g7N;F/R,1?+_G-ePL>.4LCS3XXL/:W7N@W&INO#cW&4R:f_
Qf9e5].#6:XB50_(@bG^IeMDM5PR;&A,_D\g==J;fHXTW3_>aWf2O(V3B/3MC98#
O-K[SS@,FCeDeC(K8UN28LHB3:g3ZSPF[3]=1:CS1bLJPg:H0Y6J>5gNU<FVEHAI
/:78K]LVF/@PQ.S6PG4_PDIV?1CI7=g#.C>,-B@W?,@gGMdY@U^)8UNK#cBYEWc<
cP\SNRgfH1>1?b-9Y9:(MB:d=gAb\_fV])Abg:6]VCDUeJL;MWFE;WQM:>@@7=Z0
VVID1Y@1K3V,:CV_g7;C+:_+>7-6c)2eZK5,&F(^;))fA#<2cJ4??O)(=SYO]ZT^
^KC4?]]GfggE=QJ>XdCCBY:@W4:d0cbW#_.)V8XJ4EH:If5U?50^JT2g==^985?X
FAU,OD:8bWSBV+8YP=3AJU2bFPAY@UUEMMB1f)LZ#K,F?CF@c/XZc&>@X?P&A(34
89f#4OMW/N_aZFQPF:\d#D7DMW6AMfT5GM0(g<71ILW:]&+]/YYcO8@S,M(bJBF7
+G/Hd_AUF;]ZTXT8?XWS1;M(/6RON8_K\/aUag<<8L5&7V3cB38SYHK](XH]-eE1
eFKQX<\fN&-SQGF<?Be4]e4T+acF0@S@C#M#g#:e)>0BOOCGU+)1E=^3[(N6NR?K
=D;)b&APYI8>)8);\@V#XIFT\],f]],QJLY+^7;GOLR+B\8QE>(8(Ib#ZM32GQ<-
CUEf,\Z>9QY5D:Pg346S,,7SL,JW+_MEc[d8:+I&:\[EQ7eW)UF7Y0&OeZ246dFe
AXPdKcI/-6^)\dYY=f@.3e-7ZQJ<e^]^ZRa.D4aCO)D;(Y8bA)G]7e81E+=0UIcg
6^NIAI<?5+MER5^@fCcCHP3R0>T7+GFg[8&@8?IU42R4fT5+#L_:^@&QQEfD.g;;
/E[UPG-S?O7FZ<:e2=#Q&8SO(P&-M_(>A+F978GE</MLBg[MCBKX4JZ\95K)>,35
Hf)+QgZF?BMY7?H;P+-;)3H1>&g&;YUEB5<,IeNF7FI\3)XB1,K(_9dBDFKIZ<Q4
\(0LXX>#H8a+#/dC>4QLA>]/54#f:T9.gG;I8?M=QfQ3>A=F\c&>+;^8,^(bbSeL
.D5K2&LZK8-T[ZZ&U@078Z8+D^)cFIA[(bd_Xf[ZF/.G;TSYVJ.H22L_[42.XA82
.84VC:B(#EXRLc&b6f,HK\W1,AcK[RHePHJ;CV>Q^&F@6N8#9RdT1R<OT_LFaU-:
>[cE,&,;bKTW65_.@40ebI]T]G.;1/\I,DCUG-gH.RI):,JEB]#D8E>Kd:IL2d;g
7>c681V;9Q@004#H0:Tf:geWYgS.XD97.NaI+B3+g=a/-2G-)YE1I0HTI]4,N9aO
@\a]WaabE.5TP#,-@3[TMR1JIC9F8<f6^CY82;E]#-(\EBZ+:SOIN/MV.E/U8I&4
AbWVQUYNDfRC;J)68:5J&_?NQ5c3/,af]SYd)VOA_[)4E=O@cJaaRWOG31f_;Za@
IQO=9;K(-F05^FdUA#:g@de(e9[(J#69(,1E\W\7K\9DaN:-Qbe3TH#Bb2=YSED>
X+QG;KD[KdE(XS46@V[5f(I6V@:BRD113:;cce2-O?DNI:eVQIKQUXO7&MOVd5++
AB\A2S8IEb6=4-IdO:)<?8UK@9<Gg3:1BV.1YbQOV\O50Z7gF+GM4)LMR3Sb5(@,
CTZ<AK005BeGG#9Z@M)<e^.-b<B&,.62@0dbM,0@6+WBNe]3ACR#>#<>ObC>KAZf
W6#HE-/IKA83XS,V]<?YYT\L\WOg-0@I,<NRS2,BK64&cZfO-H^&.6H)M2RXLdgI
>cD&JKA,2#7=0M[dZHW?2\SgGe+c-GNLY7S@RMWF;>6af6M^]^L\<Ve67fL7^Ne;
\#YH@T.=^/-IV^<T<_\Cb^A.&E63\1)<OK&5:f<X:aQ:c;R4#836acD3KKK#>JcC
gHIWF]^7KLg,?^g2Y162J2?V/SHO,.[Pd\;-XW^N63O]\&:N<DW??U_Q&_V1.9I?
P#SX9EOKVP>,9[&;K\P^1]8,1\>Xge_U[dX;SbCQ(](gD#Rf^^#]#(:HEI=1Q].F
E9+1CH]ZJ\,a]N/32(>PJ9/?a]831KggZ7BZ6TA_a1]G^;4)PLOZ\8)2f2&L76\8
;EObY=[ga7DV#\;O6BPUH[;]DHV+g6/78]\M2]OE4.<_X#O^7FJ<I43J[\XP&G3/
fO-KL4ec0DV?^QXZE4GP=Q76V0)&7:/cgdeP(beL?Y#gHIUVQJ(L/EJH5EZXdD/\
0GT=KeEP>4TTGB^J#L64gCI+:7P2S+((<VI7Y]VI4:IZP1fD#(BfOJKa<QWS1/(f
9&5A(IGZI7&;;D4@1^7I:FNIDa[@:9E:U(,-FV:2NK](J.3T)c)>^-BVb\N@^@OL
d19^TKa8+V<,^_E_BA5JU8.ACf:e:ggS?,V^B-b0DP^UOBLYIW&AC/>(FJ^]+.IS
f:N(0<4I_L4T6EPc)FN;d>LYPgR]G,QGCEM@]=.a@RcYa7D(]K^7_J=a]\X:O4WH
TA;0(_K(1MVdXa>9(5H3H]\#A8/_/=a6Q;R9[]]^A[?<E8<N36)ON0Eg(-2,0>C,
YR.Nd,;4WC5IM,Zc0@HfG:BEP5Nb7I6[)K,U10D,N+Z.?WUcb(/#dPVDI9FO0)@X
U1[5=,Q5][4e<J?KX37Z?==N)ABabc6NS87^dW6#KJdI8b&LWQ1GUY#dbYX(a^9f
3:[(B7;LBY.K@cIP5/.DR>L;5ZEW60=e(]JO3_<;(>)CTOQ2Se7SF_9/TOI:>L^e
_C/=cWKF25TPKWK2dFSf1QVDG0I@KP?ZV(7X1&P/^RK@R-\S]b,R6e8a@VFc7@I<
V@=4/8d=+f2EG(fcR=RY@e:HE7IPKNS-O4\=Ug359-PI1>[HMdF]1ISH[H[(1A\=
+Pe28g_JK5=E,\3ODJ+NW/453FGaA8#aY.U5#35:MbDce2a^O5CH/2^S^PDP11<V
J3[OcfUfF\P=J/^64,Z;?<29_C+,HW:@]^[ZP8Jb5gH_(ZGOe[X]@?(S.?dc7d&A
^UNF0@Fb6CK&X(1f6G@Dc)@#=+7e^H7;7+)A3<&cSW?38K-&0JF<49-3QW#)<6G)
4<\:[H4+)c\3g(.L3+E^[\N\GEW#V,;>OcEOS4WW>.)X@[e#<8@Mg5/C5Q3T(0#E
W(VEJGCB&VG,+IR,Uf#+Y4,Q9:OQ@UgQKSRc>EdQ>3cCf,W1Z3bX(bO^1Td.Z2KO
3ECd3MKAf-@dR;4CfG=DO#6ZJBS3F7&5\8YF>VP]YM8U5/2I]3G>LXbCO->>CgfW
LK[=>@4gFRU>;HO),:1SKe7A)fRLc&A1Q#H[_T;A\8-Z.Sc@VA/+-N5HSdZ?8=-N
/X(_#b8RC2<c=7;BS5PYIA9YEVKYZ=KHS6VU9,KSYJP\A<-[PQ?RYYW\I4=+P;\D
A9YP=F27)7RB-FZFFA4c+::&d:68U4Ea)N)>CBVU[C=N3eP?/KT7R511A=^)ZSQb
^@:N-\QGFd;XH>(3Q-RVQ@023,TU,:\B8U?ZZE_Y^(RT^,WU1fVEM,FU+be:5D#;
bgM5NI#aba-D9ONe_,L(gN-gJQ(DJU+1[:WJcBeLP?/I,cXa(a7L.&W[aS;@A@7F
RTN&A0B(5ROX3e3-=Fb@X/8eOBO4We8DE3>1\R7ebDB)QC_1F>WG;@(Ce5IY1AS,
3ND?[dADM3Z@-8Nc[AWUe1C:g1(+Ga^3/>GFV1.=ac[R7XIF)E_9S[0\47E,-=RX
N/[1ES.Y:&KBVE4aedY#-N.POcQT-F3B3EJ:]I)R79CDGGV[)IHX\^\N>]+.b8Za
)R1&O]0R.Y16N._8EER\8JdC<J]BP^T(g7eRd/\Ae3A:M,L]:R/_/fGPWMCIRB\c
P<;58.9MZQ5eI=3SIaG(5XY&O\,]7Q#3(eWR>WaOV.d?AO@SY[3:/Z6cF9=#88OF
a^#(U:E3GTcaZO,7DGOOK7NB0,f2T,9:dbF&JF.cP2Z2KEUOQa/OUI-c>&]N;B])
[DeH,B+)SA5Y_+cSILD4cO53.dPWS:W:cQF4D=d<@c0H(G[Y][YeA1WGG+041fUb
V<L9T+D1&bJ)U9)8&[\W67A3A0A?9PbI-c8R4B=:PLFKD)VdNA6=H9ER40cLV1C5
IMYQd_&3/L8+0)/#cQ^-e=5)F/3S@D#eS2NfZCOR8gMPUUPF&G\eDI6=@I&c?C8@
WZ):\d7.FD7c])R#YYQ+O@(O&d4?AK@(N@3OTBbd?FNYES=3a-&89#2Y5#EDA>&Q
#\BR=@-K2ZABLM/f,3ef6/SU#,738Z&BNf#J-LR4-g<IR73d1<OB\7H3KAC77E20
\:/Q#fZIAJRd#KZN0d&M-8D/&XcXCV)L^=5<##^ZZB/X=&c--#0#9)Q2^ECL:)UT
.,>)@XCK#18]:FCC8]/;17TZd.HF-(8)1;)3R#Z>.OTLgBXSU>&KEMb2M8J#Dg+Y
b/TLFL1IS7g0#Y:6M+OaPbAeKT&<_6AQ919TLB^6<J2Yb4AZ>)f:([7TTY+W6D77
)C6E;P,+Q=e/3PRHU823/OM@>O8GX]SMA>3#T0]>IS9W53C(KWBB[HW)3HD[1Q0,
C>4Z:(D5WYP@XTJ[GZ2?88JI5=f7dYC^2ZT,?O?&/#/G_@\K>:FNVPW273A6>;H6
c4@H[aZgR:5R6Nf8G:J<R=AGe6[,59SfW<]US[SWb7#H-NHM\L6H]U&gWA/fbPWa
J#4AU76C8,GNOR<dF)9]FG=DD6=NFSeRg+7^[@,:8,E(]Y^>7d<9aPN#]#b/_)VU
3#gRC=042a_45VR-dQ#?aKd/;O6C\:[(12PbLK]SfcRVKV#Af6HQDT;@6gMe:I+8
K/5Q;<9bM0IHPXW12,@:_SVB^^WXEc)P9@#=S8);;-.WNa&Z0FfIIJ\=bN4OAL&?
aW2SS7\=4O)YeS:ZQ4HGJeaG7<B^GHWFN4DDK@XB69-A1OWN?3J>8PVKJ2;F]8d8
1Y0(5LA&8MeTDA5+IC)O3OT)dBCKJ]AVc_??8bgZO<g/I>50MU#8G=G/D9ffNF\G
AaW2B3Z8Y<Ve]N5H6C_5/P9DR4W@YYESGO^a-c7(Z]X+bSV_V=;#YcF-A5&JG?4.
-YdF;33[VPX/^2F\RLFS)b,;6Tdg4+5697D(?>...1gG-X@\;8_@YD-d10e#.>9J
Fb6J:NEd<;4Nd=_57Wa72:;RIQMFQS[&P175R+.gZS_D2:A(3D0Yae&>,6.b9G9=
\&6T0:Me7BZ,9Uf8/AS7T<.MAR7>RdS+UB5L[g6C7?<(^M1+0517:&-.[9VM#KgA
DfE03c(TPf&d;-+1(bE.U+C>9:6=]VK?^P0PU6FTVEe.f<4\]6A&b<^ee<#O>4-]
U#.IMX(R-L?5N5(L?BDK(cHJ26e1>@\fOUe&EFW3Z)O7G5S,EIHK<+@CfGg^AgId
NK=_LW]+,[ARA@MSdAFHd7cE=8EJ_bN))S(>]YPK7[J]\V.N?)J[OJ/a^<+Og7R5
S3JO9M4#KR@Y5)-c\d-YCKee]?=d^A8_.(aE+9ZZ,KL^;=25WI#IDb)0OH]8E?+X
[J2fRfO#;K3&9A>[J9_)A_JA?TG<[5W-ZATY.JR\ZA.5>>&DK_WEF=A_4],Kd0PE
(PaKY#P(>)-:1c^O__4TMN0=&eP[HBX->4J2@+a3CDcHL#g.Y]<YgfYY/=[HGX_G
V&g2@&.F24-WM@2[&<B&)M+#aE@(BW@;M\=PLa3)UP4SaNE1Wg:T=>P08#g7KFLL
776e@<J3^Y^WddZ_bFg130SW/^LN9?:2N@DE&gLQB^Zc9&fN[U4[-OTUaIUe#d64
>L98:+?1L)ccL^6F3fHT)6?5@/,cXTWc#-bBbK\.Y2Q>7/I3L3RJTS5a4O^\X<EB
\2bT=V5BDdJ[Za1HQ^#2O(/I;+(Vd.(.6RCJ&48A07eIB&7ZO&Z^P_.\_Q<>^ef#
:ZU@^P3=cC>,N^eeZ98;(Y>M[_TG6\88Y(4Pd.ZWQM_+8-E9R<&AI>5K/XcZVYEb
P_SU:]QC@8U4^;<SXAF^g-9eYQ2F:<P,FSfRCN54Ef4,7c]0/]]S8I#[)7]<^:XR
3B]&EHU6?E0^8XT>>K>]X6A)/:ON\VYf&@PYVE4:2,<J;H>X&=ORa/ODNXJXRKSI
EVNZ]f^93W;REUX2\G,49GBCfCab,CBa\dFIXPX=O^1(P=de-NO0&B;GF4;Zg)-J
V_9U)B3E?L7+CDHD/UT^BcE_g8-T85?4RDSY[?6Aef1NP?-^g=-Id),7?QA]deH(
1-&/=4419>/gg?+>L\c<f;#/TY(6FV41Ng4YC8;Z5:2VNF8-;b+:@f&4]=2CdC#)
Q]1&9A<cIC&D3A,MHe6<;LB.ACO/>D?Wda&>D#Ug7EKD4Y^c6+.M>4=6\6]cFJ[N
.)]-eA@H5>_H:1W_0^^QZ>f>\f<.ba_3WW\VJ#IFa/,;CI=;@^G.T_R_c55&bf.U
Z8.(NMAEf574D0=>]TGHQRP>6<d0aJ(#ga9?&--^B7?Q5TW0?F1gcQ.^O<^_-XP/
ffQB.XV&3dJ1YV2TRJ-;_b7fO-B6NNDN80)/facOJB[M-ee(F+C[&DBQ#^Jc?E37
#7g1VH7#-.)P,:1F-f]0<?8M=1G2@cKd3-559&GL=;E&^_RWOH0cO5.F:I+L)#82
G(<b7^RN_e@[BX69gc)0Bfe_M[G8\e5-0K7WA?N5G6\18AQ--X###-VQ5XAJ_c#Q
O#GXB:TO2QA(\)b;>#M(R[DN4N66A,]cR38Q_5;V[dH_2T6RSZD?Lf#P#:?//@De
592/f<BTA]UF-5N9DSCM;JX:C)<g-J.YH&Q8S7S)f&<S02UABDZRD;=9DRUE5(?d
]<B//;;3P,U>(FSYWE-ZK9gSHUB-BVb@ERYc;3e954ZHIZfG.c;]^c^OJbM0-^]C
.1d.bONOdJ,F3\\@C&fSOd@.U&6H#></SE3&QE6RY,WKL]LgcN>cY^E_X<;)X+&1
b(MeK8eB\-)(N<)O_.99KHZ_)VZ)<:GaJX-cH=S/.Ha0:;[[#0-W(_&AMQ4#2]a;
)U>+eFWNM=Z;3QbB\a/A:TAe0XX_2)@E7YT&4ZQ+7TGeFgHLC,+WDDIY/E2TO#?<
2WOTJDWA40S]#?:JJ])eBfFJB@e&;#TK8f?EJP(3-FCg/;,EU?(g,_>TE#D#(I<T
f_68^]W?U.L9\_=O9U@aH;8DD./AG4(RUdC-5W0PgKISO6#MfR;,##B<14(K-#K?
<W(7-3T@11A/Sf4=XbSM^:I&9Pe91LOHMF/JGcQVLS<7IBHF14;@d4Cb+;K-Q-LW
:F??<8Y]d<=_/5_=/bgMBT@M(>=YKB#OTNH#^QIWaYea&9(CWPS@70)T0FeU3dd:
;G6#3N,:<>A_N[SKR_(.@(NY6_#VY)AW>4eRdQ2<J_IgFNQYYICKD550g./N-FT1
?U]VE8R_Q&S7?&L]R#T;(R>EH07MW;ERcE:Me;AXS(AMOeWb9LZ0PYZ07XO6KN2A
CNB+dBOHRQ7B/[+Ta+A84]CM@SCJKRcT.H]JA2HDaAJ0c3aa\-[?d^QWDCF4M]cf
?^-Q>GKZYALUW#5NZbVMV=HMB6O/0]D6TE8AUX:D,)#K>V1&,.+GX+AWIX,K09VJ
cX0GO\IG0#&K\?&=XEKMcN6=<2I+D_[-X<08&MV3)?[KY@86_Qf[:_BRRY21L-IB
96R=WFf,Y#?2;XfAH2X.eICE7b+8IE.G47G2E<dU.Z_WV>a2E3:Qa9<##TV7FO8<
NFaW@Q)BZf:ZSZG#\WVDa-Re^-WX30BTX4@;<gc\dK^c,6gOH^:IZZ/1&b.bE<S-
-3N_,d9V?aJ,aXF@S7cU(AD^-2WXCB4//YgZJc)7Wg>1K:+7CU<5ZK^/H1bJc8Z&
P#75)^H9,:)R&CMU_>P6QGd4]32VFJQf=,Mc;/-=D4O^OGgMU4[M?&7IID7RN@IJ
dD6(PJ9Ec&O7T,I&\=WK)HfZ6RX+P(1H+FMR^0fMK5+U/7#b)5aXU4V&#)=dYD[8
9?>.5WU:J#Y.9\JI5&,V(#.@[WY[V6I-[.D2(9;K_:OJ.@-Y;0IE&2Q#I;E>\<)4
=ZJ6++01N--cE[1<PVe)5J=cfaTZ-2Y:eN1:.RGICHQ?)07Id4c3=E[^V=T3C&LC
HdJLG9^F61)\Z^2A?HUEUc:10-:@U^^AW6)VPN-\)RG9ZQY&USS;3-]VVTJQO,@C
9M]aRY/HJ8&PQ>3b1aJU8CeBK73[J8J(NNe.+YGGO-L=e1\.0=Z\H#,NM/OE9e^O
FIYe438b63^c5+d1#P+>WK9_XfU<2JOK/H1BL8(6+^a6CV#R<.a5#@N7QV9-GWN&
OZ2FK)H#aLERRVX_XR:gc4U8\==Z\AAa#<c8:P4:YgJ;1\7/V-D&;#?6<#\,]:Yc
O(NJ9JS,M67/T3H>;4]S<VIK67cJBUfIR1XR7Y1bN[Z(S.N7M9Y[O5^e1Z3U.9TK
L8bCYK[,QL^DATeVF?d286ZRQ+&>(4b+@SZ+b&fR7dT+NB5]J)HK<?V(KRbSFfG+
D0V;4W]Bg;0>TA:2W:V&f,+&^Y&DDc,8RRV-4R&f\#K_\+IfG;YW.bWf6S-QRf]]
(WS8O1>bG#K<BV&73a>:#<HX=P:aEKO=(O96@I&<841V_0Ic]AQW0Ze9-Yd#d7L[
9U[1AU>BRF[=.P6M?J8&@FT5[-\-O=?_5XZHP-g8>9FK-;&P0OEgT)HScU/3?I_/
-Q(K#&fM[6.^?L/VBU0Va35CJ;2.^7@XMC:PN5[8eH]DgcEDM@4=>1NW>D6_D0f[
SWf[/,IDSCL.TBa6=CY(FTZ-I5Y6f,J8SOH;KBN3De]VKVS:6^;fQ>OOYZB]72C^
CL,aZ>a40P_#Z,1(YU^HfT#.J-Te=efH75+V6Y<=@>M28LS.QC],3/.J^J\YR77f
7Z>E4(6e57TcaLCGZX_;G\#5A4ZCR4#??0+G.Z0;B/c=_Q)(;8Z_WV?^-;N?MK#,
RCU&cY&Q>TdF)Tg^dDI@+>gg5-6._Nf@QgP)F<H<ODe:I6@D1N2(b+WebX@XB1XA
FP.@3TbWUF=C]V#_9^eb=J5^B9f8ARV_MgDB47+a_[TX9P/,DQ/V4fYNg[G6\0TG
J\ARQd(3<OFW\WTC:)N7.G(-7IdM>,/R:I;L,NfDSF=8>/RBd8&Rb)YS.TegDLJN
5=1QZC;=CAHXY+_&-&.KP6,H8QBBXB.6/d7T0O,V:WO@5:]D_beed7A/?L1]C<Qd
4_YTBPfg;cA\.KZD-ZRMOAQcTSMV&]0+,Cf[f(;[N#\4Zfe4_;^b&=_,3<JI6-a\
^fJf1.?O?2IN/B>)8HJ,1/N205[\B&bE[9:?(SZ[LdQ1U1.YX/e:^?1^SM-T\^L?
TN^9:J>=BE&:.7G))g7-2YB0=TV5a1V44?-0X=Pg,L5\@+;,F73M/+=S()T06R)X
2[A=K1E<>I?&8Zg;5aPQOJRDUT5UJVdbc>?#-+/:B-_0P[Ha@,d80FJ,\FUYL&cV
?4WRfBMJ3EA#bVf:I-b86T83+gA<&C/^HC-3;HR]I:JUS;ad@\f[J<0=(IIK4DQ6
J5a)R<F,Q]50W/g8beRfG^L3J:K:HTf=O#,:VOOgW.HOZGa6.Y?LW=N1c1S>=5=/
V#Ng6F:C5&3\F;d7fUB?V7I#T]:FWRN9A,FbADc&0GGL)N24g-gAUF6?SZ^3KG9<
&]<]]2S#0dW=gZ=.\XdgYF/J2e)C?NXWBD5637-[6.WSK3.CaF:>3/ZNOM7L]7Me
/+MNfdN79Eg40NVLTLbHQ/B#87B4@W70:ZQGX1@,#<UR.>Vb\KI[8&e\5#F@@7g;
(^[PSRD@,F#=W#BS)ZK6V4A-&,Q)bJO:9?ME_2C)d)U?X@./e/&#AYb+U&:1\8(4
7O:=J#W4N2BFGaOC2O>R-3LYN_Y<<0+WgJMcSA10\3<WZJHaK5W52U?N;J?S1:d]
WQ3393V5;aRT7S3XFIeC8IX;26T6+?Rbf41Gaf3J?e?FC<^N]>_+EG[&O8RHZ)(A
EA,g)1T^D2,52d<d>+N#T0RRS6@B34)Xa7EB9XF-GA5&<:&#ML;A3JBdV7KAM74.
X5&.JN7d4GBZBd07K8R7e6^LNSc>(V\)9cXV)KeL/H]A^UB]_+2AEEf6XGGZ/(L_
;cdWg+LB/EG8#H>HOQ,c[1(bc&0\U4+4(7,+Jd&Wb&3bTOLKM4#fEaIW_@a^TE7W
:)IMHNbHXS9]\C7)F?1\K.PD6)^.V@cP((]cbP1N>0&c]FbMET-<+^4N3Rb.^I41
LW9E=^#dQ:R3CX._\d4_FD+,OH;_)8<EgM20:\N._Q7Je@2]/<W3fQU[9XK/0af0
<W=bVMaT0R_S+U8Qg44:2OUES.0cZGO4d&;BPO.7]1XHg(NV1J/bJKg]:g)J[&42
OJ.g0_c\]P;O+DG#+J:2Q<RXLIL:>#Y3]248G2W&IQL2^+QY]?]fe[3DW/G)ZWD?
^M#+7I1Ja_+:Af<U#cN_0U\RQ85MX\7=<cZ37OO.I#C1^^&fHc#D&^=4fd\>dUS3
4STfZNfU6DQ@BHHH#.K_(IL4F&9fL_VcUF4+2F^/#0R7#D9@KLMARL/gPXF^58W-
+L6Da<&U@##6P0B\@YQ:-FQ(GW@?SH7&:]REJ3EWa35BP+[QaKL<,K;?LE9F]1]T
g.UQT</5bS2D._AZDZ2LED4MG=4OUV0<],)M<AHGda<0FG?W2a>X]b_bMa6+YR66
/W,Ie=7D7)@Rc\42_,=8[\19O?:DZGWU5SIg^P)MgLS,fH9UP1fU(-4/VW2U29P\
4ZcgVCZ+g5?.L66fD+WZ;f;.+^^B2#O;/VV&5=,]IBZeBY2Rba_g_VIbaP5.5R@e
,cQJP1^8>-&D+bP1cX2O5PT@QHM_DO5-#O2()21BBA\CAIe48QBO9BLOe#&4@5QU
3>.Fa;/-QI>3Pf-KB^;>_VKV3M=?g01fO)45E^3R]UR3=;EBQ;0cP4cJb5=Wg[H(
Q/I#/G,PO=1AKTUC8I>,_TALJS\;Af-RYeF.=-.X1[Ib22XM&Z\8A>;L/SP==601
f,a@R0)-RO5Z=@;+\a=^gbR=F(/W\<Cc:91WLeKcU/g^d4QXW0)7e1Y/.OA@^>^C
,Z]5Y7\#0,JfHR4K_eHXP8T_a4N>FQ4^6Hg12Qf_4G5,X-#c&O(6JG-Y_^NL+5c?
>0A<&I8cA1IFELLY]0+1#I4>HRe.^c?3JCTAQ:DZ@+@N]D3#F#gED8U0B9YGYN[6
6US;32]M[).-/7@Ja>bR9Z,P^3P<RSL63#E72\/2<2]7Y[ZNIHQf>(d;,I^?1T2J
&.F2=a+I;SWOZfbLV)Z@[/AfbY?9]4?6,1c#V(&+3HMLbcDB<TbE:2>/)M<Qd^@M
fZ\D5e3LOb\LD83CfdZ@B7KZ/EC(+aMMV??cMZ?1>b3\f-^G2?aPOPCH_]JQ/2d#
gL-PD+9@4M]O0@:^N_RJ//>?MW&U&BT>W;ZWdc+,dF]W7+Y,](KOb_Z,^<@X7[&V
-eTX1)QO3YWE<^8#LY8:X5EIPAUT3_=_RIOWGH(EO2OZFV&-?F=&40TSQ)eZ?M;0
:.4]K9D=2g])I?C^,06GgQ&-V,D\U_FbNF#0KXP]]=.f5OJZ\#\LPBSGBG7.S2&?
:f;T&2MHC.=_F@@:HgIW[@)(24C@c2O/,P<O4S4FAG)5]1,DG^2gS/6++\G>.KY<
MfeB.FR8OOO&YSM_>+TYY&A+7Kg]X<HNL\\G?2KCX<^<YRCdGS@&JG6[&;YJZPK7
->;>#]1g907Q9LN5X^O1Q=g;@/f7IJdJ)+3YJKWYcLaQb1I9L6adCVFT[)_G7H^Z
/ZO_.6\R-?I=II5M/(g@HF5e^MfF9-g8XSGU\\C<R#5&BDD),+<>Q,__H>XE4.a&
6^c&J5/cf;AHBUg2>+7?>4STgQQ>AMGPRRGW7D^2(]&/H6D#6]\>\eP8#330[(D&
.H>YWeEc8f(Ga<;^e_JeQDAD(](@Gg5Rb4@X/&FTDV>VC4#c4(DT9.cG^;SCCBA>
f#=#Y:QSJ@/=C5:Z\&2\MBg-J)eFEQacW9BK9G7I(Q,a9U3X@X7?/-/.6?#X7@dH
_\Q7615YW_AeSNc)]ef,R7=NFX?XMc,5F5W+#35:Rg2/7e,;fT:?ZYHfYb;BJ2TP
aF/K/agdQY\95K-/6A=,R496RS-YCJDLN-,P8RLgA6B_D+R/1+HaV;=A:S768J(R
9<5WeTF31Q[8-T-ff0>S=#V?UNR#3dFb2(U)dA+Ea+JNGMQf)KY#::Q\1N1Y)Wg/
C[]T8EaS(P[(V>E0)FY838[7/0@/7BaW/4[+GC1#+:+aTG^@,3KDV3CN:GMdD4EM
T4;RGU042:#)S3IUJ[1c#d/.&KQP6M_Z3=N?UP16H#^=8+72W?KP[ggKGF>>X:8g
B,U5FKP@Y/B/SCAOb?5#GX:\B/P@.ec^\HGeG/PWHX/X.2aKa09V/;c]ZcD0Z+Z+
U7];Sg2(V:NZ^PTU=QP:[D+(?d4]Q4D>+8IC[DGZ:7E6+TXSL@G#2:aH/K2Y?<5_
.=1ebc^[9KfX-MO\dB()I(\0,e8XgCEWZ2GY<-::5R/Pb,BX6V7_<@IgdC/;0AV:
GYXMRG4J9da=_T0QF;KRBVTW/&aaE88.#SEg\/aFF9.[9C.d^DS>XTabX>9)UJJd
5GN.bLVX+W?Y0J&-[YCaN#_)OJS>?,PJLKVdTE.G_QL_XS)Nd>GV\g#C&BZ/+]GF
_c\[G9+7UV\[LMK:4#+_UG1R=>YAYLDJXfK1]6+WIU:8\(,F^)4ILfgcL.EZ^>K2
T4f1g3JaNUPe7a+U3ec02IW+@[>4E^04G8M0,fPL)aA&2P823bI_=+MPJNLJ,<:C
.CTL)>b@Y#BPT^HY<8L[;=\GF[MLdW2[-cDHRJU.(/C;RGUZbVdeaFH\VXS&Qg0G
(?cfYIWPV6QOdGM]f4W_QV5-JF[W^6H,X;c4JE/f-62B\5^NC3FVW/<-S<fU7Q/(
LI42DP<S-4f^_>BV>8fRe&VLF\H]05?Y6a8MWN\&4bcB5(-VMc,e?M08(c20_0b]
dWS2V;\S;b[UL1C__2g8Y>EQAGKH.)e8OO=S)eG4-9\E?16(CI.X^\\c\98K)0XD
MPW>HME8^Q^fDP7<3@a)5<S7gCY<(0CXE4e[-L6#5MKB;/21E=#XLf/G(WPVR.R/
3?K>Dc49H8<9/0KTgV\PGJ@+LPS7]9HE\&F5gBg7_&L2d0S5F2:<a75^TDSU2fCJ
?OPL4>FFN.)A6?W>P]CX?0[5C#@;]d;[=28ZWYe:OMHgg7=H.O4;Ue[Z/c+R4+U8
,]GUOHK)^]3I((53HIdWc+2-/)YOZ3^?EQ..dC.EM>^f_B<6C<F&E+PNffWPO(b3
a5.8He5+PZ5[Jf7e>a>\c?-DE(Y96d[7f&a+1,@,gO/?:YD_0Q;IXM^3EWBO9Z\Q
OA^&Y8N4<#3\(c41WW-GG26Z]L=6422,D\-V;GKG)_>-IXZgMEYP9W:MZC72\Z7Y
+XQ8<JZAL(Y6\YSeHBgR.9\^A<G/G9=9IMgGZagCPS@UFVLEG)0/W6IF3:JYE3T-
PYPF@@V8_SB>69-X/:>\Zfe7\G-PdP[NG9S89MNB4NK8?EJTY6gN6\2[E9</BNeF
ICC^TX[@9gUG9>FUS6Dc6NHV?GW:^]c(<dPdZMT()>Ua>S.VLSHQ0+Ta,a&FTV:J
]7:(RGO1Hd>a+5QK[5Df3BZ:Qf8#OJ67)(:KP/Gg2af0S&P-EcXY?/4E?6e2JANA
g+)SL<5fTSbNf0[87VcVbP98Ag7>JCEN;B.2,g/&:ZIH=\>74E/L69UI&CJBZ]bW
3gG-bST>1bEZ08(1VG?Kf08a2977+?ZML(L[+D3>=9\3+FNB7.I]f_[IF58Wab^4
NQE_5<M_6FeO=O6B:;P(0MH:A5aeNR5H>YI)[,;K_+AWON9:PWY479QQF8;\eXdb
PQ@?b#6O2Q)]TL>W83,\I3&C3S-E,)C1_#>2e\S[KZf.IOAgZNRfSc)YZYGCeG#<
?FX:K?;T-GbD23_-W(=^\_HdOX,<MI3a?RR(B.+=dJ_f9EDacCP<AP6N:T,b/bC?
OI\C9X>&)/:YY(@#)[O6SHf17^9_4LF._fL&GW4<89W<be-=35[:eP\J/8KbDMYM
d;/e;cE8e8/BQTSAY:f6KeS5fYE(A+568S+ICPC>f]a\BQE^8FAa1/\T^7(P>6Ge
gA4W2IaXcLbND@\fI\2J=@JUQOD[4-##:eLJBLg0U[/DA-e?7aV,G^_,:\/(P8?a
YW/G@)cH\];[<_YK/B3+fLV5OfW[I#M+c5FVAFKA+?@7CDPCVVFSVRa:3cHQF8J:
e9(1[D#VSF.>O+T(T.8K4d?c+#+6Na0TUdBPd+_#KZDE&2gKV<8Kg/0V1<9-[A0W
DP9;5:X8eLK55CgI:fUXF.W/R+AaSRNG3N7-CXd<[d.=QEJ+D,[MLYcC-TRHLfXL
1480Kc\cA\.K=g:E2O/YIH,EdNOJ2\2P@^03E7d./13eM_<2-V)ILQcR.FIR[+27
G0db<2\_)),\RbOY#4WNDf,8f[G0R?U&6A-Yg@65B.g5K?=D_-d?+0T4QVFfPbbV
KFU43X/2N1(_JCc#LJLL:QMM=P\[@98E4:\&J7DXXAUFd.#?YQ2&9T_W/34I06Ne
c.SRZV)Y60LBX8KI&E@fK<NCg&@X:8:#8-DF_W.aK(EfaQ+bL>+#F,1,bSDQN8)8
N<C>MQ@F?)K&J4EASHfeR^Fd?H_Wc-CW.&GbH0OQA]@F6NMKHG<^V<EQ#bCe-Y@e
<OWF@6Ybg4g/4OZ#^IDQOE0V-&TN[[g;<I7BGH-)c81JGYGc-:5XM^+V>S#<P^;6
<e_Rd/06:,U)U26)WHJ^[.XC7+X,[C<LZH:[a13EB\8b:5WH=LQ=:YMC>#H]Pb.I
FXb0IZP\9g9D?XYS/K0b\P^Z)5BNZOC[[R-\DGP&EVQO_GI=3cPe&P8^<cdK4[/4
aTNY>.[.V(AWIc>+CNG&fZcUZAMV5X/XCC7R1403>?#Q#:YL@&5VfC:bHVZ6Q-OC
E4,5dA\dBU::;-.fO<JCBI#^GGDO2f7be[]=7Eb9J/dY2+_>f]=]0<^Yb?KWeJ@4
SEZNd8(-aC^C<<FP44K?D)aFW\a8c83S^D8;LWN7H2JAXD\(-N(GISWa9E-UgUJ>
5E31OC]ABJ/Eg1.Cg8&4V];6+A.^<3g.^Z#9RE/G25P4L4J[2;#BG.42XVdFZ,/0
3^6BRaX_4NTdc>-,fD8GVe2AHE7U#/+A2I7?E_-bF+C,26@F?SD#V.^d#IFULZ)5
E340H7:BY;#fcEPVO1?Ld&Z8bF#32>[G-ITdge/[Z7&<8JXEf_6=f]0aa3aN<Kd]
@)OG,DL(5de-29I/FF.d-5JSS=V.YWNQ^\OU8#-,TbIH9b\g2G/NVN@_YA)OU2_N
YLa(LS\SRQIE=Q&]1=LU<B,-^Y\7JG-/[1&:NZP9J^cEFU4EN:X=URDORG(9]<]Z
\fV#O&.<M][f;Lc@M#Y5cY,3=6:MXO@O0NE_4Z)U?D9H^F_cFU@W8)BMa>ZA]B84
IDT3E1?&F@7.d>R/OL,A)6=(04]N=9JDFgW2.1K]Qb_NB)M@<H=POL>9I=f&VS-Z
J0\:Y&beRO^[@4HH8HLDQcFQ?1_\fOdg4OL:?F)@[:VG8=U_deDW57AEZ^@IPaaE
GU[YNNK[f9#2/PaP8a)7OY1NV#?V13II=;PZd-\9[7CSMHd\1:PZ-2U@?6Z<Q8_0
O)+NHK>=GP5ff2a8V;=<04RPI1VHN-64_)Z-I+96>GLJ8ePN[BUBM;5U1T]HEP]M
^X\)[5D?.SJC(2KS8XO3eL5TK_Sa.SD+53>QVA&GJ@@&OF>X@BdAXNAWI^b,)E\d
b&>#M;P<<+_S/7]^:0SKHNdY\J<G@Q,JGJ9L]fgV)&S^I#8+L]YK89E]aOW)H-?-
A6Y9XA@D9Cf^AQ>@=XGNUeI:<88T;d=cV<]RC99X5bE@?5CW\.FUX6@K-)>Dd9=S
5<ONK,EfM0&P:d.I1ASbQ]_3dSQV</8NGWIME1>;Y1W,2a/@T,G66(]\KD.V8La0
;A5e+d\KFFN>/IU:E,(NZVgRE06WTTF>5:RR,UU(G91+B&C.RQf)b)QF4(BR<:/1
Y\MHT4@Mb[F2dMOe:BA33E[,RP:OU,IW+;N7a3J,a,I^Wf_A]^;LN^N=c6-HF@J:
]UVaI8(Y<D.#TCU+bJL-E73ZO(,9G/f=dF/OD5BJ?#YXU^D/g.W/e:f=VcO=I3WU
4AF?8YRV(Z-OH<\a^gWaTLZ/If<A@Cd^>fK@g<EJZ/)b#8+A=<Hf\&45YMW#d)(X
S:4(JM.PW1bR#_F/We830a5S69e0\+M^+9)WQaI=De_)JWf=Z=T&3,4(A:Z>XYZ?
<C-5+DfDK]^R_IY2\d5RCFH9g]Q>AM=5V3R=P]F)(V4ET9>SQZ6cBV4X_cRVaE11
TL([=Yf),dX_cc/J>6^-Pb,/7K8,;<7&[b=XQcJR=.G^&aMC7]4B?c)4W[?Y\FG(
=dEdR7RV8C2)SBVTS/N-LB(QE>,KA[d5\]bYe98F/VBD>F4>=VJHc#Sc1@>^\UWR
V69Z_F=S-E.^.W1PI]c<G#LR/)M7X+2d]Z&8#6H0AEDHNP=-)MCf>C8(9\62^^0A
2.RYJgb/9+X8\4T[CM(Y>MK^eBR_g=?)T1UKEKIDDOV-XE\<(IM)RR;eR[L^.f3@
2]VJ08,cQ3XZT(Z\G2QP>E5E<b[U2TMc(@g9G,bK[OM<5gJ&<(WY#]Je<HQ:bPKZ
A@JD]A;_bDg8g(dP_2_DP^?X[.>UMR@QRcdKE5IXHG&-6867e_d2eBDgAUTD6;G0
]d9D\N9Qgb+M(;IaSK5K:3I327HJN/g9L,MTD;&Q-c_4Z-[[.N]cd:LTfI::;dTI
.Q/X;/_2#NADeMUeA.:fSbe4-KQ6ZPb^QJ.3>9KQ)9<gKMfQJB_W=8[cYP=)NfM+
.c=.5.I5)J&bY)PLb:BXHc()<Rf=Z9EHA+g;55GGTb1(a?#/dRYF:BSYGQ)>3J)^
P64>7bBKC5<Q)C[0\+8)_-8d&1gZGTgJOWWE0^SB76b92P>FA\P;3W^PNcce3JZc
:CDJJOT16FgfY/_^,?B&?/#>5J)?0-\>OKS7B7cUcWf]E\VM6/H0\@]]cB:?7>HB
U=c.#G[BdEZY2F_CZ]<]NXZ2_O-d;.LA=--&D=,aYH<cVDE6:^ML4L,GO,;2cB[O
@V4)c;9,gS/J&H4H3>_P?EW/RJMVaG@O:A@4S^;MK##&HV0+8D^BQE;V#T#XHIa4
2QJE+?X6R^9?+V0-=_&/gCONZX8XM7[.V<GU_RYU=U3WLc;1Z6<;ZN>f;Da,7Gc3
bWEb1aDUV(#4X@[8F]ZVGB<KRPW-YfPB2^F8_/fc+3I,O?e9,KCBYRFCTE-L5+0O
+d\?7E4UX7+H&9Rd_YU&[FY8/5Gdc1SVK-AK?U:]CddX]cJc5L2d-BRZ49],1BdI
b:R<;^gQ-(7V?,<)R46#(+9YJ053ef-PBU]KZ;eabP#)<8b2/^Xg=,@M#.DZT-_G
_SK36A#_\b(WHXV9\GB5^OZ2cU1G8#3T_C;WR,/9LL56-&XJN+IZ)3bWO#6=2[E<
TK^L?SW/.OJ4PK9>.PeDJ1W[-GU3.K7;+-/XW^OPcXb3VX535^;(LUTG))]Gf/M0
b#<DQ]3WM+,RC^:PS,_U^0U](6[#RaM_MH&ML?H-OKMHZTW=NcYK5>Z;LY/D#>JC
QGFTgJWTI9=eM2K6@U^764I@_E:2]WRA_E\NeSYKGT_3(/=LC+1fK6PCM)gDWA5V
\&3=/f;<\VaIX[()5]XCS\^X.OAE6aJaL:T_MH/P^RB=FW>cAH[(=6QF+.H3]I8Z
P,^)TK_4\C<(N@>IQ7P-aYBR6_U@U9dB/6O@=T]D)@eWHO905Zd-OT6fUaG;(T&R
7Z81b4K8](@cD^<N?O@X5KHS(]#7K:UY20cRF/g.5=6#d50OL<aP@;,1./.-a0\V
4=58U,]@;+QTS;,=6CcR-^Ddc[=>4+<Kf7&F=8W6^ZZ#[f+=9=;@P#RcT^\:QN>&
8]_)3Y->@d0>G5aY@Oa>>0SXgD-eA62#@^11]]V3=dX<3N2J5)2#.E-^X.)E#[#J
(E_dPK&:KU06Wgb4dEIVI9T)FT4bZQ>]+H47b7V+B#ZUR=1VJZL)0DJ#)[41Zb;V
@:6^I;Lg/1R@GAA<;]CJU[Dc5C_Z].6?0=eI_#P:Rd:61ZbUfH=/CGa=DK[H4a8;
:E@O6-6fFK,H4808IE3Q+>BO4X:bP7]2K>92=A4DWKY#F;K1_2>2=aL=QADR90#D
E8ZVWXZJEBOB3dA4M/G]J/8c=75?X;2G&a-VFHb1HTPT_]KK0)K<\=[SEU^WH+g^
3;.@d_83:YIL@M<(Lb2K\_(+=4FUNg7e5O&0Vd-gb8FA668dX>C_XF9>UQg:/e=L
-+\@XZag&)G\U@=>MJNI=E0:;:OB^cGJT@[Jd9_@U;:FGJ5b->NG.DD]AU#(T9H\
PSK^IH,C=K)SW-6Qc3_Ge4_RS&#)QK;ZW9+g3S3MT:cDL7[4=;g=gS([[.S29f<:
V\W^BeN1XFcbBVdcdM@\AV]L)HA:Re^4R:b,.M=:K4P^Y[5fbcHO#_KH9J8c]KGV
_2-MDZBTP[Q/[34fFaTPOY@?c-IX5R@fa2C3?F#=<7:d+bXCOS^J/_F]C+2/9J0D
#.gT#BeQ1=2[Me[Cf/IRJ:]f.5=XEaC&,H^INJFU21Z9-=+Fe11MNSM-XSTCeRDE
AbCNDTgRgVU;g[5bZ8X,>:aJ_84(5:0#SN]^GVM+=cD7JA<93S2>c?CBZ-^_CS_?
N\,(<T/E-#g07G.LFRVUQFAAY9eI.U^JcO29Z<\\dIHdf,[aYN^>dF#gL^d9J(LO
\UVJ78B?4ZLTgd@?D[V.VT2_WfWUFZ==>Z99d4cMKD<TZM1cdg@]>DJ,MV(G\7f]
1U3V4eKRLI,7)QbdX:[[7V07-Qdb>)#>9E&N2N<+K.+CX><?fUKO+23CA;J^GYKZ
L^H]I0EB:O7eU^G@P>X_1E8YLb0?-O.]+F@RA@H9fYXTT6KBcSKPc38b0I2].eVR
BeCZC#cLgB<DU?.5\(41+gR97DQS:?U4gM[@HZRY=R6WGGW0@.5-^ecC01Ta^\PM
Y<gZN,<ST(K)#;U2fD,,]I4@#CJNH#=POVfNEB5A]9=A6e,gbO:P_5UKF62f]G)e
d56KAeU/[GDO2:FG@_?4/K6ZW?Yg8Fge^=^W2]c?N?&2(#B#cL58BQeAY[UgMZeO
Q^:JJ-/5>GA@OUSeW\Pde>_A<+Q[ZM(BRHKA1US=(K3O6YK81LG=IA=]OF0R_\/R
XP_,D4G0LXbJEUF]<=]2_:OTJU(_,XY0+\JXcDT_H=GMIe:<S/F>a5=,1J65@0N?
^UWAFcAM0#N2.Y@cBJ8DQUS_AMZ:E,=(Bc&K&GR(4eg_1L78R.[IT8Od96Q#39TQ
#DE@,SQKDJK^>)MA6JV.J4aH:08V2:,E-6g,X@g_3_4K2NMY]9Xb.KRI>=]LG\;:
cJZ6/TE<6Q_BQIGS9<a3@;,_@M;:ECN1O:+^#3W.gO6K=]O;d<LBZVIO:Jgdcf<,
0O1W@]9gR:4Y<dG^4^1E_20L4BV:VefBDY/5ZHR@]fS180@^A9.4e>^]\U;X\>3K
+BfT37@HJWDUM^gKA8@]W-H0HaIN7_&:#L7/@8^&@64>S.>\aE,_2I.Q_^0WGRa@
XLE3bI7Z0Fb/JU;9LZLM9dCJW6X278[3Ye,#5f3J0/^e)e]=K.,cBVb-eJ.Ng&>a
L-[_FIZf3SDOZ]@J6T0VDKREFK7&AgB<.T6]Y)[_g0DbL?-K[8&8I6_&BGfU;A,:
B2E#NcV)(Q,?aAGFg777[1A4c:e\a9PMNeY[03M<+XDEPPf;70)g8@-4ALOJPb37
Y0OU:?XQ@If8I<TZ4P/BW.#7OPb8/PTG4PQ;Q55)a8:>.J=NZZDTbO,/f5@^d6#Z
QVGZQc0.cHT1TX0#V#I:;=<X8DB=2d_X]7;65#1)#,1Tg-LWg84Qb?XF\L3gHJP.
@3JD1EJ7+(Ra+?Ua1176XSP4b92]_Ua#_/6:WVa?fI=820eIO3K9)H&UCF@Xa,[I
O.HV]S/LFAA.g@NO4SJ4=^:\F2Pg&aBf/6IA\[G6&_)3\>SDAVW+,_L[XYNOeA.(
1V2;O8UE<RRZda]X?8T=0GBV1>Sga+YA?DDCP(XVJ6:DA(VU0F7((Q)PYSK7NT]K
KN6(3bO9,RW,P:2b6TB\V;eL[?P1\,eg5QW@I^,F;D8R5RZXJ&bf/IdeBCV8@1._
053YZZG?.d6M91e0FLC&YH<;bK/7U+I],O>OJ0:,L^HK;=S_)=I[7I/[GB:YVec-
LMJ=[gJa,J9eF;OA\D/H@BFdKYG?G2[,J_HBSS,,e)BDDK1R<d82T2UF(JC6,gc5
2LgJbL_6b]A=dSeaP@H&S.90P?-SdGcGMaaH\+<<ZX5#?RND/U\I:BdIJS])U,+/
OA-2W5@KU74>Q1g2SaU<OCEHHK#M)X<YgVWACeJDF78YfdgZV5V)0c#WQUgBNN(7
Y,@Ifa_C#7.-_2^@2db-9HY)eVBPTRWHR2d2+TL)@OQM3c08?ObP[80-]3?/d,5f
W=XV:#3gH/2CD/TK+ESIFWAJe,Vg&=_fcT@#VCIBF;A]W?1Y&T.Vg>,G-Ka).U=[
R@^G.JQZ.A8C93\^_=0<#Y[9(+IVG+f;6I:OH3g24&E,eDe7[a&U[DDgO7V<75d1
;_+f4[U,9)CI9=b2;XFg\^(UV>a5-PfPK0H:bI27ADJG99>RZ3<,T6_?/>b:WLA7
g/B0@O:bU=[\C/S)gZ&@IR8I^R>ET@FUL.-]17ND<+SMV5dG@2LPLV0aG8QVCg1D
VXOUX4f+\W&-/BQab0(MPM)3ADG^UN5SD[=5:aH&_-Q89U:7Y(B5M_=_ZTTDLaE,
>K4)@0Ad;_Z_a#4f4b=d64cC>S9)[:73PD48<B24W+F#:G1WR_R6H1gI]9+/Sa+S
Ueb-Q^[;I89JDQSAL)HJQ<dN&@1:_.KM4Db2;Q1-/:WD(Dac<)eYd.J9=\M[L:FO
FG+=+;7)5E(bb,a?A0#A+fc9SJaTU;M225C@JK>bA0K9J1:eP<YL5>^]U:>B2g.P
fH0#P4)WUD\8bg\)fFe\BJXYG33U@Q5D)>OZ#UF)=5&I(c+a,Z1bDY\]F<2FPcNf
E;ISFPcPAUK<fDg&?9=0AXC;5))VL=VIQ[#7U1cGD96X)I5E>+a/R<#AM>:8]#Z4
Sf._VG+:AD1JA=[>I7,AMdDEUUY_3ZID4f3ef59:I49GNc_Fd,f-OEB0K+/1Y^(O
,dQ&RD(@<TMG:ME1#S1).9T,8UDZ:8=AK]XU4C)b+APM+NdYWL9YFK?Z/KEeU=[>
B[:/BSY9_P:[9Xe4]4U=EI1T.X#)4B^cf^C.L3YdYe&FdD_X9]]/eH25GHf7eD]O
[Y=2V(6(>7#3gdWgK0M5aegDTW+LD8CUTD>QOgA)/,^fD:SVNgK^3W,[ZdA\KZA3
#;c0LN([JNHU;RF<Z8c@\)=ECRLSUJRC<(7O1@[G)7^+a8M]P0Y=XJT-P)/0KQd]
M2^LJ:#U\L/NB#(Q-LJ6A<.J.(Wd(>_4W9R2Z&=PQS-@&WZ/X7:b4;&9>M,KBEA3
AAHH<G;;@KH0=W6+77_QPC]F:7M).E;X3Q?.L8fc4?/XA+^R;bd30HM,DJdDT>ab
:.FK98[CL4_g;72T:Q2-U@8]T.CGX\(A>.+B\WK9C0^?@:<44E6G,3@gaRT^gX[/
^M-O7B0NM,46QK>aD\&.f(3Q2a@=)O4<R.G]3Ja?Wa6C/3XV85+T56,72(CP:\+[
@@_^F/SBe49eeY&73NK:NBEQ)<C]?)ReJ6BBVQCG/JL]gRbTT,_8^-<gDHIb#HM)
ZB^(\L_?[8d8U/a6Y:V.Y:T)WSHKVHgTF@YE]BaU[O;Ye[MBE6WX>^b1Fgb5^5Td
X>>#+gITg?:d,U=2\,9HWWP=[c]X8caa^ae5R7?aH,4/dJBN3\b[fg/?ZMM<?a3:
Y:G&8@+TdD+OGKTK6.&7FG0@LQ1T(Fd)fK/0SeY\@Q,bKH\gD)<P/dMf&S4U^E:5
HRG[GRLO,aQ@W,/^GNd=cTf4F-aaJ?R;&TUfKQ?a5F(#G[_Q\MgGILTb^FTOAX[9
F7Q;CB;LgQ3EQgS#d8J4-GEgCK89:L[=.P@0U>T+@-#D6YW7B&=I]eBXI]a-OI7,
?[\POG9T]X<UTJOS2(U]?]<.4LUO4bca_-N0X6WW>c/<9GALY5U/;dQF?g+YX.,E
cSDH7M=B#>O=B_:S&J?>M.=IgA&.5(T-LL;0Gc0a9f(5,2I9.:9U;c.7;Qf>3a=(
DX@3/E/-bU:6&>8/KG9O>;#==N=GegUU8#[\J4@0/D3Md.M3IN00\C3NcNWLB;>8
K0Ma<LccbP=5)CK9N2g^XU;F-Y:S)Q&32fb,CcNQBFZ\;aUV405(QUB;&X85+gFI
YR[V;gDAYS@JdNRZ\aV<7B]EH>J:a9-_19?C30<8BN-FMd[#WX?D@5=FX]7V&DB2
AM?:Q.A?0_@AU0+&Y:H/O^Z@2R\VY\Y6X>3\P(0L)R>.IK,58K7O^=W(:-+NcC-\
Q1TX^D9#99LMQ-@F.0E]AU>SSgO(Y?26;a#QGZ3Nb86ZJ;);83f=6e&^A_IN4JRP
a5Z&8NEDH7]-WL>42dHe^.87C(dV#A)C_XT=G=F1/)+7:SPIb-_,(MWD/=3O3Z6I
W^F5Abd8?PB^=;K=cQ:C<1?:d@K]a?P)]?g4CXg7]^(aE7)TbBZD47GDZS7eMI[.
Ef_[]M,0Y&-;0(9.gU:N9)O_LMHJdLG=Ra_U=Tggf=_1W&4]QI+H(GLIc.RNN2_S
I-F>TTF7?_9)IKLF,U]+7BT:.UMZ^K+#NE+;KKU6SJI^UcA()OYKce+Ef+dIgF;6
gSZ8[><(M<#E:UJD8]82:&b/6O#gI<K0#:>WCLD=>IXd2QN>=JY/e5(20LC?H]Wb
W5QMV<L7^+C#A8d;+L\.SbZ=BY7G.eZ<VF00P<J[]HSE8R;M//Cg-B##eRZTddZW
H:^.8EKN0M)-/TFe<Abb:=\)05=(/M3H(-2dQeT7,8b]3B+3P,7)_I_cO^-[)geO
?_R4<<M&H;;d9(J?&U:@C1d<#WML\U]]aQU.KDVB6T-H/.K4/<4=Q5UO^gdF4be<
]bL0(:6KU()LcZ@dC@J7d);B3E?JW1T1^55SH&16>3U+ISI(3CIRJ/,,<?aI&CcA
R#RK;PGTd+I-,;KG34P#<41.2NL;&e2&LS;>7d#Y9Q^WVUJXC[SS_7X(a<NYLPgV
W_6WNPSfGNK[5(]Q6gV[IMOW=e>-,&N>V(OJC\9JN:,GL/H5.NKG;DFg=<VaV6STU$
`endprotected
endmodule

