`define CYCLE_TIME      9.0
`define SEED_NUMBER     321
`define PATTERN_NUMBER 100

module PATTERN(
     //Output Port
    clk,
    rst_n,
    in_valid,
    in_valid2,
    matrix_size,
    matrix,
    matrix_idx,
    mode,

    //Input Port
    out_valid,
    out_value
    );


`protected
2Pg@A9gWdEOJ?H+cZW\c9Eea@JY:-#CS3[MJ?4C-(Z7^MQM_(D)(-)+&9S[]HM8Z
c+NZKNNV.8=T0ZfEIF@OH72DW@OUI(cDfLAOE<YfM0N2gW-UL\Mg_,,K,.\;f^5^
-BfA+7=WW8:a1VJ<ABU^7=95f:Eg(4R+U--8aY[EA8,PK((N/]#2fNa@LP3\,BO:
V,:a&HI]E7Ka53]SHg@]b;N-.:(8COXd,TK\,Y#f,Ib1d_VY-6TBW_YdEU3A4X+.
PJ^9T]YK=eL[9S;QS;bT=@=^)L#M(e73+^G2f-]J5Wa#6Tc]A^=eg0YdK$
`endprotected
output          clk, rst_n, in_valid, in_valid2;
output  [ 7:0]  matrix;
output reg      mode;
output reg [ 1:0]  matrix_size;
output reg [ 3:0]  matrix_idx;
input           out_valid;
input           out_value;


`protected
N,2V;54YQ,NJ8eOe\&@B/@.3bQ;V[P+Y.SVKPH:[:9a^.f3f+d^]5)_5H5aMUN7R
NIW\e];AGUcA75>=7d8C(4BAe&KLgY.5ae.4#@;_:WgIfZEgQ8AfJC:F5,WE^5SZ
CA\N.RE&&0NQ^89[XQg0eB[@^W8gHEdL8__9+bW:R)QZEV<PA(+fZS,E?c&>>;-.
7#\_Z4<>9HcZc,0+/&:=/BRA:e+9bK@/1G[/RN;@[TN9ROM;5]4bR-1e4dE1R9bJ
SK=NfA,GJ:U\Fc).3TRSDAeO/T?1.N0X)1U+R@ZGHXS)#N;]6F.b>]VMc;C=<a>L
9V1XaVM+>S?R4P<B0(:cTPQF5eae&U,SHVVXNJ58[eJZ/LK-_U=H@4Q:FR\D&6(T
bC7.f?7YDPDL&#f&X>,8<F;5@_?OX9F\:AM^<RHbXc3aE]4=Mb]&0GMLW2a1cE+J
GVa?A9)A:&?LF:Ye\gJ7:>aW9C3=XVVT-X=-::STOF7>XdV:;&K:@&]]ARP-+/eU
:AccACb.WfO=9d3E@G452cf3_0Db2RF@CXW\Ag=bLIWd35TIfU&3J+fa,/C.aM#S
A3&e3f2#D&R[c.+>;^g.KRU;Ca7Z4O&(Md\^aS>>JI?(:T4fb2FSHU;D<[J+a+]@
B01-9/f8;LH6_?^G>I_aP)^GJPK[[=\6.5/12A4Z]C8Pf9S=aB-_F7U4=N<-DHI@
[=AFS.0/DTUO\AVBV5+D&\b7AN=Fd[8CRC)bOSM((b=5]4@2[SPA3X;C/-+1#E-^
&A1.BMGaF=e]Y?74cROgTYIV:e@ATA[H7CfP)6=?cB8U+fFbSKNG1MHb<a(+MC4g
S@;[B\ES(AL#C>C&O,NC,Wc:LB)OPX1CJP.\874:[5(OLabNGMR^.gS;cHb;2\eM
8Ha?eYWWHca:06_O2cLBA3=.P0(/@+]#gHOC<9;1=>=c5LTB-/B1SI0(W>#O_3Z9
6:52/5=b@#ELGS8fZW2X1.?YA)/YPg?9+0J,&TR>[IF;:>,^Fe,K34ED9N;^FFX-
BC.)MM@/@01WFRU.L-,g=V3K\Z3^6IGe5EB1X3fV5QE.Y@CacbOf6cCY<@DK,#Ke
=IV/8>&;eD@.=>Y&YYbDX7KYEf)SDTGZU6afY&.fWZ-JKb\MLP8UQ8QSQFK&^;a_
Z+&N,4IPD?FOEdDO?\7<M5S0,?2ea_,83gO<_0GSW/L<.H-Y+2]Y-<a>e#0;LWEV
K(0N^6L+\4_\2[GH;b>>R0aJ1+UPQ#eV/^\)R6Y^#g,KP(XBfNSZgCdVJJNg#++F
S5S&aTL?YgWOeM/T5AHZ^6B^?&DUP)U;\M/1S2Q:a8X1HMXY\4Z[]I7?=.O]B+<P
:[/I.fD4UB?XCC9861&F\g[YYeQY8d^-cdB=WACbN@9O[;1Wa[LVB<H.;E#de4Q^
L9]FTJCVWHR4Z0#XR<eHYV@ZWH_b9S.6EJNT_;CgW6b3H5dVgJAdP6gf:[+Cfb1K
KWYcO5Q;OL,RV0gIAYEd,LP,JZdQ+NR^/D+;23QI>\AfBI4bLNMM8)FBP>9D-T1T
UaX_&egC=DbU&bP@R8WD#N)F<.^QQVJFMb:@98)3U1RNO](D33N=?28?O-#J.e#-
([HL;6,EXDULP>;[C#<6V=\bBDMg)?M)GC>C328,]#(LdI1DBE,GHG_a2Ug_)G<<
CdRFATDTF#c3?.]1^,]]O]4@IQL?K;C6BZ<,\#@F+(dIF99GF(5Ee5/?L:Db91-N
WN:\-NQ177gXPaK,eXAfN=ZC9eV&?U@X=0I[4/S>^-T4AVQ0QRTJVD3Lc\>11I&=
.V\6Zd0ZYS+@\-0U6eI>,3SN;R5Z=5C(gU[1NXb4dU2?VQFA?T=(Q-Z_T#CDM]YV
/@bQc=8)(a7KO?G)7S.K_Ue_SGQ4R:2T/KD<#PO?&(WN9AB5S_A,?a1B1F^.@Q5^
)YfU4D1]U@I82_N=cg1]Z@:]^]a9T^fQMc=OYaKPTU;N>Q]QBGU,fgM\5X;NcbdB
--Zf1O.Cf7[P]ZaEM\BObP@K7E6OPAOa;?PLK^D+\=(Lg>]IR^^DKV61-INU9.O.
3<<eC^3>+YE:7;G0@7:S^H.<-_9VK91eO.+ZVWKUJ]H,d2WS#0,0DO6#f9]1\E5P
E5IS#AK0R3g?=LZ:1Bd9<=K:9BQ&bMQPZXE7E[#:JZdb>Oe,5/QSB_6f2<-90(K(
0CU]Hd@R-g0OaHgV#)5I[caNT6B,7A_NbGPaLZ5\PCIT=MFNEY^E;5C/fB+3c:J:
<@JS/6T2;3GK+FUHS^K6(PU(V6O(@;>LB6Qd9?>LI3=N1FKOI&]=CTN[<&TKd,FM
2F5UVDZ2+:_/^UCB9W+,RPYBWDNB<93=#Q7=N73A7Ze3/:gIcKgf.X-5\e<9&332
Y\(MS3H,R,I^JWSG\Pg35D)aP5dP<eE&ccHV3;QMZGcQMO:bJ?54a.WWDM^&+d^?
a7=\ES4JY)\XMdb=<A59>Z])1BW[];J&7T6P-Y3:\0M@&FY<=RD.U:J[ObQ>Hd;7
e9R#]ce1>-K_<b2R@5<9I\.WZC\=JTb34XODX-CIUU=0E#Z\EN85<fab=@8VO-80
@K,#1&;#\@f;1P1373b-;aE1-@Y\6TO;<VW446Zb&QYZ/A[/0?TGWc/#gNJ:+I=/
DXaEC./NIdW_gP\MZI]>+2aK/5G?FBI<-K17II&f@PIS0:SBD27OLLEWI5?J9OdI
0HW309d]G-UP]Ag>JDAY=5F^BUQb<35E,c29H\a^5.ZGPF[22PM_MYP6Zg1:;8Z8
7GYVU.K4;9.K49T[U80BCRW0+G_Z&,d[dWM@b4DA2/=>52AW8NH<gDLVe8&Y95X_
[Z@=,LV(>;L=]aY#/#0CJ37MRAR6_;()gE]19BHA(0<?O?TYM4\(L^-BPa#UOY)W
aOH;GOD8?9^L:;)agYGGa_=]PBE+V2D#Z96Z\;d)[7PXLX=Le@.C;DN<+?7/]0ZW
D</7T4+&KYT2D3+U&3Ke@>NX,AA)M+?4MfP,(:GJDS?NcFa]@BKaIE6D)gE2P>Na
_9,4\Kg3gBBEfV-8A98^f7DdP6eIO<DbP.Z2JaSdM;;f?E6(12W9gJ7(DV;5a7ED
;-W_E<&Ra+:dQKBO(fAgO:Dc+B.Y,_P()K\1b03X09949)PGCdLg-F&G1,Y,cMb0
1>;HD00:]-QZ;9cYNdfS.F=1#^AZ/#J:T#R,Pd,6RLeaR1FQ&daU59S5D\/0WOFe
AL,b:g+P[Gb]07He3Lb:7P:X+S^,)J#<Z90V;<CSS,g&7cS(,FY=d:HGE<AG-Z>#
AQ-O3C@c]9[&-R)eb:,)1cYM60]XG/d5_NV#-BdL3CR<K@[:fG:K>>3D/CE^4e<5
6GEWDMU=.C1@LZ2cXJ=bL35JNeQ-6H[4>a4\7WUACJXK57XS</^OFXT+]QN+[;V]
#TZ)N,2-fg3\-9H9=/V_T+=<g60]gU-/2/@@SUED20N^d&E=WU<Kae8_,^4]Z8DE
-Agf7F(AC<deE)7ON)G/#(c:aKNO,2ed,-<6Z--,SC^MLI2,\0+F.4J(.&0-b_6N
BZZa1F,B=B,:<I[6K<N?99MV5YY2732IAV@RQ#>R:_-:RJ+;BC6\;.-ZAJC6O8gW
fM2Pc4X6BB1@E&7O4Z]ID:D]&c6V99DgK:Y#7,I8;b9JARR+C\Gd+F#M(8fWH_SD
1Xgg37;2_?+g=([_\^a\9a[0W7^DP[@1FV;S,XT/0NHSNFJ/L(a]=>\JK7Z\YXZN
;;P9(@L]96?2=HAYfCCG8]#X3VV7>(VB5/:fSX65BUHF?KcS4IEK<U1GMd#+BTfH
/LF1HL.E_9/O8V@:+4(;b(R:+-f6</VW\9BV_>5NLZf/1G=J.,Qa6/T&Q](8+HU-
TI.fB?_J-Fa-FK5K]A7#B7N&C/JO40I3?I00Z3Y8W#^WQBgXP0[OXP]26=&N).WY
_+GOE&(4a2;8P<f-_[7aA5)@.29IR5IgY1?9G;XP42Z5P7RGB4)(_<;Y7CfEGI>c
^/UG?AO9^HX/2W^A(]MS/P4\S&c]#X5:ed5\Lbb4(Q5W<)V^FI_U3aLQ):MJfg>\
7.YUVDBKI67K/IZT[GcLN\:?QJ[[TN-AN>]HMD+9A06U+1VHJ_Mfa#8/86K8/D]&
/2,WA?0O[[Y/NF1U3R6@MKF38EdLZT9UX:#2Z+J9&F\[2Yb89<P,gDe:8V;e3MPa
aM]\/?F,8^5AJ#C+8eYA#\HZM-I(A0be+Y(YJ::eXS>\X7&a6<S1V&aM62[D8dVR
23(.V(LW;&MSEbCX@1P;ORJC@U#/Yd?MUa8]2FN>LY]NZG7438&ELNJQ6FN:#H;d
4>#BB&.6J\KK3Sc4<?J#8QN^DHDLZYL]0^TZ:&9KPN@f/B_F&D90@:G\S42e__Xa
\_4TXU;Kg@T\;&0[-NQ^2Z#>JdT66EX)f0U8Ae4&ACE)gYN05KB(]C:Z\X0g2AD9
QFNV]41+-BWC)C0U4W)_,?Y0T0+KXa^KJS.db24ODTWP>:gZ<dB)c]UdFRZZf)ZK
5,<89=f\a/^a=(XbOa8a@cBd<2\-2BAcXU8W@+9K0cB15)AB,RBT^QE\>=:C&g+d
^Zb+cT:LW\2:#2J88XKU5D3(0MDMUb,T5,dN)G0Z@B5.EC\:;D9OU;@b44)G7-Ia
2C5@:=M:#-\gC5Vg((9Yf[LMK>97&TSH91Uc)b1HKa5QJEP0LK6S]?<>G9##6NN3
gZ[dC/&-BW8IY(9F.a;8ZUK3,.NU<AAERaJbIAaf<G0eE>DOUCU9@(dGf\EJa519
E+I]Bd@-fWYDA1M.0<4UTD@-\Rf=L?PQ03[]8PHZH[UeF6@SR<,?.?);4IZK&(X+
,YNVVI0;Z.ULZEa[FEA+YA9/6Ha9@@J76Te-X]EQ:-M[7Tac8.7[2T=K9cd-4@>b
W;eJ-2E.X]<6_&[&[,14VQVOPQ:McM)&bV0AXW@L/-?83ZK.#,QS1caL]&B/FRX0
<fO[,a2#Q_8?1PC#B;_DCRMbHIcGUWDf](.FC(/N+/e7H^J7#=UGFfRa1NaL^+87
<,&R4IgAE-XN&I#R96^F?=_Pf/W(3?HaOM>HT_^:Mga[.gBS,0\G06&;/?><M8LI
-He4#f2KO.4FRg(db25,0a8E#=+0b><T;\3S<(63-6gCNG-2g1E@FVIN_]8\<>]c
=)<-^,D.ePMaCXKF0#8.>X,6#2L@XZU/fK93^e#aL,Fe,-_0LLUO/OYf-5VS--d:
ZC-[=Q#PI]-Q&ELJ8LCX)6fX]C+OFX2ETB9)69+?_DRU_+>2;AERc:97dKH_WJ]W
bNV+DH+=FUH=b-Sa]bG#6-5F#eR5(>daH(+C7/)G/OK@7]Q8b]J9+b_\(N1HKdY2
AR5)&9bE5&gF2[F4&^adP20#O.M[Oc517L@]W.LV.N;BY?P^[J73P[@(N9fRFI<O
]d4C-B3R#eYX)<&I09Y83XXA#BIfCX0?J^[GcbP>2.7^:Z-\GC@E_:(&0W>,=KMT
/=TF3Y_:7<MN?bEPe+5ZNgAf&21F]C6JCf]0gcC2^;]Se2(]QVcFg]\<;CB2^:F\
f#)W?[&K&0N(Kg[fGgRY__CX.@]+GcFR4X99fL/ge1WDG\<(:;JG5I/RU+Dc>\dg
?0,<4X(FK5NS3WE)dY&9c+fb.2QFH-2@CGC9S)b_PP5<Od++c8:<FdG+O+ceBTGE
<cb;62B1SU,BM<QbaOPc9d6#e^VHD)/GcXMT8b5.Cg>Z-gD&gWdL_fJBCQaM]]L^
DM2KO,fQ@ce9EDYD<O_LUQ_I4S^MBM2_DeTD49Y_&30-60TM>TT.>9a5H0JSW>Pe
0>..A@J+7CKK+5c)VQ1;]8cVb@6LV\RO3Q6/8?FH+a+P3U&2_cdd1+/7&&?N,#@U
-(+@,ELT(;]<cHZYf=E@,Cd1c#OC<V3FL<8PXBg0g</\Q(<C79^73MD#WVGWAbMG
?Ge7>E2MN5U?>#d^2)^W=D@f.XVTS8.B>Z@PI/#>_f#=(Y+7O;\@dGH0+;9U2&SR
<?f]B5YQ.aLB?Pba68f:D)/YKU/+9F-I?aN.::d+(;d<Fc^8;E3/9MfRVZM.aD,_
[f+7aU8KSJ\[=.FV58+0D8Z&LY(E85b#Y^dOegMJ<VX&0FF1c6XPJKI(<e1TO\_B
#c:G<F]XIYBOcg0,7=/YA[K=T4<1Q3JTES&dD^(@:GD=b;?.f+aReNT6+B>J1I7_
E>H<YQ#F=96b-B2TEM+9^PKG5Ng:(]QOOFfWUE1@S])D#Ce^gZ(PYD#6FV2V7HA/
]B[Z5UKUccQU2EbF1/(_FYG[E,&^I&Y#B+^6baNa^Td/X_cFU+dP@M/5_3L&\#]?
GfFae0SgLWF2^;9POJ?/b3U:C1?35Af>=^O==f>[Z;;E@A0NQZ(,]1B?/)2(D<g<
,F@SLPETaF_\>IdF>>J@?HP<RB&]-<>+-N,WaBfFXE.UP_@Q17eS<bDX)^c4V\=9
;5D94cNg&V+8U=bG1GeDB;FH4g/K3_XX8?<V/Q.<,XbA1KWUEAGQJCW@P2KNH]Bg
[Y<H,V8<U)gM4cPY?S3:a]fEOBLT8?]SUWgS4]E1B/5?a<a3_-__/0\K/1ZN2SPg
P/3+M6TEbRK8OO3/+YGSQEJIIDe_&]QQ5TIC>.-02=?>-TCS/XQIN6U9GBNCd]/>
9X9B3<6JQ9W4<fdLRIeK-\MZg7W;b?6<NT:]c,[3V#OAc0#d#,G6)\JYT\_=MbdJ
BZAeKRZJZHM9,Xb0[A,+eNYEE<5>L<S7D#^COB[6_+JRW^J.KN.(3cPR&&BfO]cQ
D_@9OWOJU,Ha:eDBb7L2&)9<0b7(6f\^B(LSZ=6C\4eBdM</^Z:-6-ZZ#R_C+Q.\
c:;L8#bB3)D]#ZcP;XA7\N69)gTEf.SeWSf3]d>Q8MW^K9J#.cDdV2^4T5?dJ:W>
Y8B+&bW,2_.8#;H?63[7&XG/ZJ+J+O\V#dI&9O)gK[=>,gJ8Q8U_bc=6B(F1aG21
DV[[V]A00.OZ@fIJEe[,@-4\GU0YJC;GcRVEG+5R7[bN61&4E)ee0ZJ5Pa:SJ9Zd
dMI:X#]bYTGYcNN9?ZZNKV[c@eF]YU(9bGHHLXUaN71SNccdE\]MQc<^/X1\(=38
<(3T.1KgM@DT\d,PFY3-0=E3?cM;:XcX]\Eb:4aBdQ\?:AON\UFa/bY:dE0,-E.a
ZR48.cA91])&O4XYe0;W.GEP49E+?XL>\3fd&7dfSGB@3^C=PV:LWML]Hd;]_X[d
dK_L3\7;g;FAd2c)5F5Wf#a_3[9]5RHB,>MW=35F-a]ZVO>9,R5O;2_0ZW+/f,HI
AUOSDTX+]/4H3O)P193H.\RaFXPWaDg48Vd[Df.^](]O.K\DHUXTf?SbQD+_Q4P>
L_>4fPJd\ZX.af@^cb(a1LTf7M#Q?B)c)+0\gcBG=.Z=c_RN_3/[ODeZ@I.KHKY;
#=6eI-^4?4)L[N00+f=J(38F6-KaSTZULH1/39Ka&G7XBSL2gSa68@;+:&_O6A8V
-0SbSX4;0@+X/<D>A7M,-41/e)_5TEWWXLaHFJ3bQOfB^51YCe5,d2T6.,I;:GS(
#,?64.OXO,<@]D[KT=/,AQE>3C)D?ZTEgJ+FPWJdU+KdJ6_EMGdC3@.dD/c6.1HZ
X6&/@A3EAg@<HCCGS^BeS2VD\KWdWZSG^U[#0dE0d<-()Te]A<VIZK=W.O6/d>]@
0e-WR6ZC6Z1RZ[QF4O))8/TSVYL+J<_R,dM7dF#V0]PWO)G./8C[();8622_M,>-
-(ZX?EEP[J&4A&Q0/#@/[WXf5:ONT#Ma)S+bZ225Q/U<;##GIDS4SH2e)4X](89^
fDCJ7XG/a9P[^dG2#?E2/+.FIRN;4RPNYeO+023QQK7NX\#^7U<ec>1<PJa6TdJ^
=1JZT\/L,.R<>=I)1]>OQ[1[YMRa^8+NA?d16<aC</TI\<cL8L^Ca,CKH>eGT1/0
0ef5@5.+\e-H8OH<Bad9^g82a8,8N5&8g7M--b(&4^GC<&gRW3\?_5-HM;5_1WYb
TdIA3>VgGS;9:HSD5Ca@c#C_eLW;-E(a_I>LM[>8P1K.0A7OHW\1BUJUcNTS>NeX
?ZAd&7J<YegY>UF=,TVBOGEaLV-RVV\B_g\TBZ8ZKe\-2bH^cV^JT]X<X?I))A;A
FNC:@],FK<7;a=(.4;>4LfV9DS(dF4HW:VK8JEK/Rg&f]V3+d3>R>_#6;Hec>LY8
V/ETU-J9g4(e]NHCF0>PN+V@#XOS1>5U?^EF/S93d2KFV#[Ea1X&VC\6+W@dDA1>
b^MMO=CCLW,O.--NVG4EV.M]G&;QaOYHDDVdY5bIANO3,FE2@RSb(8TZ@OK@?8T<
&?X^cSVWQ7=6<QB+ba,X\1@RGLJ,+JTPL9bU[^)CSJ]cETC\]W7K#4&TS,=If^N[
bdW-AF4/>D+XV:X\CSN>58H/>fQWJRc[Z#gXNR_ac0NgVP#,fS_V4.5]FVbGU&JG
23[H)YNODJRf/,H/TQATZbSMa@6dG-NU?9</cg4[;NbEcX#WJ[H/Pe,_KWS,T](2
H>>2CdIL;CH=7FJ^,Fc5/I/PO^X&_:IZ\)C22XP=OIVf6E-,dZa;N[#;c<4VWMV8
:G3;E_;CC/BW>^_/O#J=X3&P7f?S0.;/?F8^#[PE[8AAG?a>U7GeAe?W8gM#2[S=
5TT6XNC-^#7G=4f?:]?V8LK,;O20e.ePB/<IWa(50.&Vf2++;e&:9\&gW44QgFW4
\8-eSWC-F(3Y;g?99Q47^QPBR/OFAQ.)+2.FL<4V<L#QL88#A=Y-P/U2TL1)I+FD
V0J(:Q.8D8S8K)3=#==B.XX3BK6ON<M&g<dNON.GS?W^WL)f_Ac;4]H8EULf&F+:
<&2>2Y.2D59d66ffHcP@:93c2cf:e5.TF(;+?:^DdO,1B1dcJ/eFVJf9SOg\WD9V
&<?&:acK/6_SN_I;_<W6H@=S+Z\JC]BFRCJgD/\RA76JKDKQM3J8RO5bXOVQKBa_
(RaEEK9?L?W10N=((J1^,RST)R_](O96>(gL+B/Q5+MNLff=#@3e.TM9e4:+83aY
/9,LK66-QP0_WHV,bgUA6bG[_@&3b]#XgB+_^DG(#,[9)[YDZ7fU/\K@>&3KF]6X
We/W<cKP>;DWF[NL<YBBW+H2=^__OdGTB-T.Ra1aE^M=S(I984WKP4P+SRdUfgC9
_b2QK[.Cg=-=U\X+WfCEcffbagYL)_CVg>H=?&F<#8)a5>AHeOW;C:^K_\&ZI\WN
9X]A,1[\@f;?#@cUFKMB+>:da>WZbD1OSg7,F6_17bLN;:.@C+43^);E<\?ae7CJ
^I>FFAb)E.Mcc^R?H_JUE=ZSV=B=]06P>)c-Q.JS]K6UP4P3E6WEW#dfO7Z0BK_X
?GQ2&ccLV\>A9)=\-<\UIVV0Te9ce2KXH)O>I5@MIKOMgQ#5_H(;QEN=WU6/cW?W
F\XABK^2M?=PJXB\Ea8H#1Z&WT\HL8S=^B7IdgUB^GH6=\@SIOGPCS=&2(GZA+V3
2bJ/TJYO6B^-]R^F&5B)N+N9GAW]LLZI4G-?:P6LG>K2VPE9),;]Y]YJE7WF(aX1
5P00=.#@G+ZEUdY/883;L]A-0KH>Y3D>bIX,TCO;U5+JR]f4EL)/TKGa;aZBQ1]e
NT]:ZEcaF;GI=N5fQ9,N&ZU;O]<<4:gTWJT-Ef<LT85Qf1@B\(Lc&)E@c<U?B^^]
ca\&O:T&(\,#U:P&CLcENLZOMV=GdX&HXSA6ZX(-f\Y7]-fRQ@])+1V:@7GA..aN
]4+6fU^Pe(]1AUbBH13^:^Q/L6YLMbe9-e<Igb5-/\Hd-XR83\X6+a\PI)K>W?,,
8CbF24HW0GDR&4DF7T@G.-=#Zd7<C2H^VD)0LgM=-R15E_._eKSdQ,;V#=:>1DHB
b&BQZV.2([Z#2DQ6G77#&VI^@X]?Z_bB:8_fa@Ed?dg/WFOYgHQ^5:N9ED&7\6N]
?NGc=F-5I>=a5O]KN+(YB2C/=WT-/fM)bOfgFR-2I@6SR[DVCfK\AV20C2@K)d?-
>5[LXOXC\RYVfYU<=DS&@(\1BJNf81XJ@OJ[=G5eRd,_1399;EV8f#PRDgAFEU_4
9CG>\gLb0?2-[.[9eLDY;#;;:dLF9d;=/(1T@WH+dUOVT3UG+ZEF7bF=DKZB8#)A
e4;_8B2([UHXE8a]+05ZTLTa,@GQ/CDg:GX5F+(D]FZ7\=7CTXE:5aJdKBX2DNH^
^A..8BJ9Y0_)bR,\=ID?<@)B\5WQaSU&S&WAeRYF[HET>B;391V+0Yb[4TUU,(4U
2@IS<2aEO;2QZ034@QD.<^[aE(2J=Je8&;>(M@F,W,U9GYNUE2+-.;g&R6QC=TX+
1XMge7)+Y>->P4.K>\)21PAWC.[g]-K-^K;AU<KLIDDCcbfR21TD#4[?@R7:^<Sa
:X>MdARK4H=@4e\SU)8W;d?>R,:H5cD1Z,867T1J\a2Pb;^8?5b;60DY-48JLJ<W
PB.?A8:&J_->+YdZHaC+d&HLMTX+SD(SW7\C+b&R@:?=I)ADZC,1^e3,L)Td))dL
,LaO>[^Tbg&O(Ag<H>Ya\+[cbe]]58R4IYQKZD4(8VV>^O21CUPDMSPgY/,DSE>g
D@X=Z_M5RY<&f7>/CC16/#WLB^_FY/=fS[Z5[.<98)10LJ,\0(ONHRXeITH^9,eY
657EF#<9(4be+J7WMQFB-PW_#(75P3&d<J5Y8^_NUgT=Q-Ga6:@@B7RY^/D)Nc&@
F[T=AebA<4e6@^Y@S[3;7)/\MF<_Q57cgS@beM5OM119Q<G&[73][d_A(;O9;GGH
@:K.<AARb,08712/,5UAY4+IFKfGLe5+J[ALbND&AQ1&@ILZ\IU)f+bX<NEEJSRZ
aD_IS#BR^]+>APP0LLSFI4;b<VE/C<?_IV1BUB9K/Z5P68>S#M0S]2,5])<VSL=H
4J^)06V)RS1:c._E.Kae^<H6:_Z33.NGS+:S6b1ZU>2g<36._)I;HU3UG.MO^/)Q
59ZV5Y;(7OH@@O=<aT4<F_eI1.B^R:Q0=YW,fZ?eE)LVP,[H-DaD_3&U-4?.B@RZ
Q@-6VO1cBZ24VYU7&07X7YKdA--b;^-fAe<AS/cZ6_2Q#M24\#Y@AF_de>7.D/LP
=)BTc6)BZDR(C;MKGLP]Vb(B.D7I/=.>OdF=[L;-.d:RMba]d[ZNJ7gMM;\ZINW.
=E8=X+/b\;g:[]OM[\);dWA_]V/D8OC/TOb1RUKE:=V.f:=QC6OR/H1AEJU@+]J+
CY7&);ZQf,/>-aQH7V-3/@6d@N-HL_S99SD\808=0>Y;2e=;gDTKO?=_<21N18]6
TK]DbbT5[P30H&Dg.RU/XQK2#Q4HT-f4GH8E:Og2P_^#(FLVaY@e@MSFVBPg_=CS
0caH3/07&1-@c2gg65F9(NC(_8[4Z,;EHW#a5AZC;JS;W2e+c#L\,W;NTeIE3B^1
B031-HVbQ,c;?SgBQ\7^)K5)HBEGU]eC&D\F<04D6G>DODOVFfI8Dc><LgEB,/Z4
eUFD:F;a[>:IKUd.K6I^1&U2B.?VL6fA4PF7.#]I#Za\C+Ia_dJ+2UgH2Fc#>XaO
9BQDM0W46-ZYgD^AQO,cPM=]5JV2e^LN9<,G8A9[85TELMHH1faW:LJgY?CJN/JM
O5Z_]+8^5IAdY49CI>VXW2=TAf5:3#+g\;J1.bLcQ))2I37NLARVZ8B_.Q4C9-2L
SVIUcD-]=b?L^^9_&(4WG.M2Z3NR<OJ6Z<YbZ?c_eYBQ<[)J^fcB]/.^bUU@BY1W
462&U]>#N\Y125YT2H[:P8D+X5:<B>gOOg+;Jd1dA_/+25>I7#]b-FQPJKO=H[__
>C]2d^U3VK,BaNV6)Q3^<^d7U:)UgH3gaWO;3J<B,^MAOUZD0SNFS[38J3aJ&f9Q
cT;L8.e-.S.,.9d+9bUa+D/3)E88;<&:\T3@(CB/>)/c&/9LPdEKZU4#0<e4(V35
)MPMKY>S13a1\VGHBf^C(<@fgM+ZJMI64.Q4&ED,P,eXC\^&A,e8=@W9N#-N3Vbf
X+E&d,g[DDNL3a?QQ92E^_X?a]\Tbc:V&fO.92/Xf_E.,-NP;<Y-?MB@/67++8]E
GgdJU0\g;a;1-@2^b^^I_W]0g0/c;EOV61N(JWLTcR2LF&<.Y0d)GCZf<NJ.=1F5
2KS5]TFNHf\PT74Le)H_[C,).?WQKIT8I@WQA6=F;>?S9Y,LUQ@><NP6g_FW+abU
HVWJE_=[AF6gDd4dNFPU<=WeC1864/RS^[:K0=/A<QV#.5,L_MT6V\T+fD07e75K
e,L=C(+MRYKc:O^eYZ,3DQW)X0@2a]7/5N[Y@>E<UT9OV#8f\KNT:\9CYSUbP))1
_ISF]R&4(=78G=L^5U8TTD2:gcL?N9AE-A)FUMMRbRZ0-/TIT-7\@J?,g_^ONIF\
,1<L?;H#V@_3C<SJfQcNgPP[3.Tf1W9_9G#E;cK1G]EWK9b1g89\.[WRD?R]+46A
f8b?XKMGg94E]R54@;7ZI)]KX^R/8PgKCA4Q;^4ZgH,N[AZB543:TTYZ\->_?fBG
H6-\8,AWM\8JA7GAe(E6]<5gR^a\OY[fQAKR>g.PI)2>^R9^cPX1a;VCRCTLL0f#
g-IZJ.BN#C@NPQ7AF>W@+6c(U=_[WWC&.c:3A4@M)29g4H:>.TXBKC9bC\LU/ZS2
MZPFRD3IY)<5U;LEc\:Ma)c7IKB+,6X@3f@5L_7NOV2KAK;W1>02/=\=1D)ZVTDC
6V)0]e1c#T2bVaHHgS\U)\@f)NNaPE4#\=<01ZW-)6-bPPg6(A.6UGPSTN@VYH=3
+@XWYR(_e=B9DfJRFL,gA&S@?&LYPTE&9&2G#3T@/aB\ZT(VRb[Be,X,b1>NC/FP
)GT.(Z7[RcQ>,3]1CL?5&XO5MXI-]+gV+cYKP,>NNF)=EKU9S=3C&J#dV?+EV2Rg
UA_@#]d@9Sg:HO427K]^J7@e@N?C?KX))(d#I#)cU_bBS7IJ^,PUW[P^THR6C6(g
Q#>)0P=L:beR8_3):B=NGHe31[)+LcI;;KCO,^YJL\=IE[\4AL+5^,INf#(J/4Q;
O6.&<O1)LSBMCX)Zd;#XI@cA:9WMP/]XN4.UX;/EJT/9VS+M?-8,K?,#XGaO,RYb
+[[JCGFLWf6Mc;&<.NFXWg=DL[(J7ff6fTYYI^7+;9HR[JTY7)fb,+N@5+F-=2_G
<-f;8a1DEX?=Y1\36L-MZUIG88BR9/#:V79f?=GA+UQO-(ZA0#TJZPdHM<>P_,^V
^)\UGCU)40#9]TO^=@Z[8d9,&^&;TO@+U9BM&E??A:+N]:?f+2=/SG9IQLADdFUS
eCDE4fRU3NHXE+6MHB=D3DBG(a8ILU+(GDVgQXW(\J,TG=4H7WVJS_-CQg0(-KJG
\4J-(>7KM&=//.]/eZ#)PT_L#)1]AF,Vfd-20@)J8>\-5X)eZ4QXcO51DY-G&B5f
)89@DKbER_KT.J0=R3B5f+90W-S:3F,?#_Q;D,)7)d^Q:26-4gSBf\&M0EH4<)eL
^?_>&F^JRFN,H09QFV(HX]ff+bC+dcZL>fCZBPJ<9GE0?Ib5IY#706S8L0d@S<^Y
+1\//<@4d9AZ);OI(eP\68K_aV)H<3-GLKGfb9U:ABQ[G4S?^VL+3?:AFH1<)9A:
7<K/#J.]bRH3@)LW>UK5+;O=8X3W)QR/4ffMFF]-?8L)\f=25c?E_GERW=[(K,J,
P.)(^:+1(D67,e9U78ffLB?dd>9DI?^C:]2c5.:XH_#,Ud//E/@>W^XOZ14_bS8>
[?c6\Q89D2=WgL.KK]LIPQ<^GRL4I0I&1H2Zd_(_6,1VF\9Z4<W?6V20D/B&):([
gUTf_L8AZ;JKgTg&^W^S91+.M1aN+f/I@/(IYe&/?8&6(K-g9/1\P)IJH@36+S5+
Fd3)B(g.GK<P<JeE+EEX-9[0A=76_R5BZH[f@GDQfQb0?f9HEHSTAR],Y=G:+XX6
9?E,D(MX9#:SNc;fPa9>KIc5G8^1\MC@B1CH8RbOg4<C)&&^AL3I/g?c=_Q9TSG3
X4J8L-C+Sc6YQ>:<P^[S_8.Mb3TfUX5P[Z:]cW2N;/bFO8MVbd:&?+J]<9AYg[&=
EN(WaS7K4LX(#_1_TBc&N;=,cSNIQ0V6g([LeLAg:AQQH29=\,c^?P3UTR+N_R/Q
2K(<__d/&3aA@<dEDI6-SeSFCP+_LgZN#VaMdH.Mg<2W@_eCHPdAS]/0T6X:U=YD
c1C5ZBX(#243I7VgQ3L@>3e]]2eE>OfV?7EIE&YR>CM6Q\RG(Ra/KRF#NBS).S6_
7[A+5(KAOaBI=.HI7eN^MXEg<]W_2Ec_>H0f8d>1M/b;cRJ#J@)+(WSTP>N22NB4
,;(LWO@<CO7c3K40Id-UJJ/_AaFeST4VEO0)OQ=H)FGT7](:NdB7Y6N=;3+e9\IN
=(e7aXIY<HBS[:CT.Jc\]M23Q\&V]:>7/H7c948PK9>OGV2FVaD4P_QRL_RdP=8>
31.E:g5:B&.E:+7fWG=E^78IHW8\_?T.[c>?W#e-L<ZZ65=30,.Pf3;ZP4<a21/J
MdAE<-JT)O;ATdC?b?^1MfObVR<(9bDLc3,P5IIeO:-S^-N6_MB2\<?FK<MRO/ML
T78(Ae_C(g^>c(#gY1KdPg]JPO]9Yca[?cPc5TX<?6<f=Tgcg61>IZA.5:XH-FRB
#S_(2:,T?=X69IE\UN[,L].RcedFG=OT8O[UBS9[T9\(RZ=f^42A:N3@\9=^?YMO
S,XJMGcRPMWQ?)K5Z=W[5WQAAQ@9P\9bd=>&Q8:=HB&_CRU2A#8>23>.5b+VZ_Na
HN:(M]YH4I&Td>VY&;G8WCP?PH[##2>8PVL(Kd?+4IT_;>+(Q5Ad:O3;0U@]QSFV
D/E8FOF9e^A^7ZNf9&=B+2bNJSaERYd.2<F)<&NSR9YXJ3E><2>QBW.cZe[Rc2.,
c93T8=f,X+_2L9L9e<4L#P_4R4D;0)CW\f<1@A4B/90/E2JS@M33K>fdRLGfHA2D
EOQFGKUQ>;[/L&O(J.=,NALTCaD0YN@6QN7QI:USJ11/B.5JVH?bTESQ;U;S#V5;
b,6^6PTW=S41bR2RaR[Y6IX&Z6Q3:;+9AQa&3Z8D31]8AcIXS.fC5dIA<UN\_e6K
3_B^ZB7T_UQIg1E@75CRHSb=\R4&9IeFZ)#0b&O>fJRLe.f&B:+e_=<5J18eS=.:
I,JER,MeHBZ#=98^BH]4(6eXWS>/<S+:@&U;-g:743J,E\g:9J8V3f1MfWMU0HA@
f[I8I0/^\0=I8S-3CK]NO6c4EX\]0+8/^#[CYKdeC7dF+<(F/YB.MV,XN/H5H-7&
?C)VX@=B:RMaYY<RdQWA;(674>&XW[W(@87C4RS9:DPWI9K/;cKN[Kd-&5ZS4>87
SR<L3KQRV,T[1>?7[WD0.KPY_.+D<9=#LK:1CT5^L-SYP</Ld-If-5D)HE6R^FeV
B4Ac&(,[EH&:-Zd)C&;e1<)RZf0BbaXHHJQ41M^)CQ/IR#L<Fb9)XYIL.J8TQRIK
55bV<P/X:S7G?Y8LZ]_96MQ?eFPYa9QN=VBRI9BJ+9d1J:N#FEU,8>#A1Ge?.=UG
E8W?O?@Q=TDS:Ff;U<(HOBPYEMHMDVBU0G:ZPM4DfC+\P7R>/eMfD77+E8M4gXD4
#Y\B<T.BVeM?J,d4KNQS+/N2A0;)/=eR>)-KfHfDOT5X(FT[2CI&LJ20E=X=3\g&
W]U/+XCQKdP0/HWg7dL7)P+UT;@D(_)e)\.A793VYCH_gX3^TUC36E0c=V<9&fA>
FNT;8;QH3+.-QIc3_5If#&[GUKTH<G-H0MP7601geYb>&UM?)[<I_CL0I1ZJc,QJ
;7aV,E2RP)ZGaYO43>3?Oc.AC:/M_R:&P07917Y_X^ZRRVX#3,P0E1Ug<,&Z,DV;
1Id(eNYQNT\@d)N2Ba:Ead)eW2\)=IGV5>_b0a<YTB1eHfEYfIL&N00PXBbHVd8U
SQ;#[)I_,fbef>A<K&VeC=J@22)>X]HM^V.GYJWD:[/UNVBFA7,#&57eT)95aF1Q
W<[a^:Y_+H+.4L@A5=#]W#S1YBP_OU6EKcX8LMQ\XC-Mb/\Uf0(#Be)S7NIWE9T]
ZEI+ad6[2Vc>dDMG]09b5?=;[@BQFddMC3&LHG;G6W6bg34RMBS?ZY=4(9JJ.6\g
VQ>GTaBO-#_e]b):))cPIa#g\FRIP1KO<1d/H(Nga^UL49+?^GW]<RMUX0P[fHW-
Wf6QX[,^^b=@L;8K_I+;[6IUS,=W]1E?\69+O/AQ<QaC575XNeTEI5-eH0SQ=?])
->?ac)KU#5OcU.=c[T^/X(RIQ/B=aZYRSJD0V>VJ&&W;35-G_3.8XR[e<(aG6ZUN
gLNW9:M2_\dKeG13a3=4de-)60LDTPSD#Ka[M0a@Zf_(G<MIZ[VGY9eR]WCPb3Qd
Q(fb9b8g-/JG#XZ16ZD8U1<KOSb#N4,;dY9[?Y)73=bX)80N,=DcVcWM2Z=C8TP?
X/9^XWIa>1f>?K.#C3T9-R31\bF:CCYG?\A;Z:8.Td/+#\\fH2A>Y+&^W(KKb:1&
R80LR<\RC\2>825>gf3bU&Z.)M_dNIR+d82WY7Z##?;dOF^\?SN;/;IQWO^P?EdB
e#(G/:J+d&Y_X]QXe9KaQUJW@[TbO:gXa3#YR[X#b3&Zf<ESAZ1YgcYKDPFM\0=Z
W,-#U8aIZb#C2AIc;Q/.5+VYCdTBPTLA::Y/C[H=-(cW6[Vf\<Sa9cBL?]Z08=dJ
3<3,@/TDOF7YMI=@8ZXPIVf0/F?,Uf,\E[I7K>gQLN]3<;/fG0[=(Z<+@QgMD#WO
cR)_D<GLgRY41c7L6b)C<3PbHg>C]e\#C_A=Ee1EST0]IBM0WY@#0(LQbY86>GHa
FIR#^U09K9\G+f]a_#:8A^?&2Ea.8_7TR>^AUHO_1Ja0[2XP[cXAPOVD)aNYY3WA
&g-8cCAd&aL90]+R_K3fJ4PZ,A[+PJePdNT3N3(=L#K-Y,a<_<>NcNPC_RC&d,>+
622g/)>4F<PW0acAR\2+(dDU4\S;<aHKb#D2[bT4.OPPfID,T_M<W:==c0/?O5GP
#7J\YQW):e);gONVAfB47#[,77:7>,FaSRMABI)eC1cQB?.?I9SPeY?>ABL>ADV.
:]bD+g(2+[7H,KNN^=g0CM,ME]BZ2:9Ceef(;&-&?A@=L;aO_(=Sg;W4\<LS[Pf&
8QPBT;7^-fcJ>[;c+SQ3g/+=WA4NT;D+)8U/82g^f7(1UgA.56(][_#@WT)<PQWE
JI1=-gbc,:](Sc,32-.P,IK.ORfPY9Z+JMB1YYUQ]fcO4^<;Y^Z[[W=^fH4fXQ=-
@6-W0#91;P,5a>5IG:QF]8Fe/g#DD?#X@VK@U7e]6J/IK(0,8K)9aU.,Z&@E&Q_&
6#MP>^J8/_KJ[#gfa@NeW,:6d#IR5<4L,Y:F<3CXW-TZe@S0_])V6&X6UI.[;V6?
(_0=.G7)HGRF6W7N4,D,D>W;PNN#K<8]HR^\;^F)f-)=CJKa:M;,:e[CQSO2@?OQ
Ff-Y6dU&AL)-#KOFT\fHD-O_Q-#Jc^afR.JYV9W>6LW\Z-Q<Q&]R]CeZ4P(]H6Qb
8AGYgT.:@JOg#<5[SS_(HWK#9(.78aGV9V0>\>0b6d3.XGPf6]V<J><HVdO05N-I
#<eKN=d>F@+c^;@+6:)D>1V&&5MX[R3]MOMZM78R;8bI0H-Vf2P=)_/QW?6c=_DP
)f:/X;^M^#-(#)G-T-bB;JA,_E?@8VG<#2@]E^/FQ72DUcXcWN=+F:b&L\MC[7ea
WJX1gHW8Q1:^GI_E4KUU(/<7@X.V?L+E=:bSgARHf>K.35-]5O94HBHJIBbU,D+e
I>)1K9be4([+0[4FXb2-_=^<QGYSW(Q5=HXLEBC1D=KcCNP50f+1E9S>b<3]N7ZL
H+HPZLd#26/gZE:688/V=?+A^H4-UGa;=,]&dU+[\4J#2<\c&U;XI4fb.1^EdbWG
Gc^9]C\4L6T(.>WP=Ye+W&+/,De-PgKOMS?D\:e:HUe]Ee0JHSOUc0?(:\8[_-E,
U@SQ]=>;Ic^N,@YHL:5:@HfNB;>aW(SGGc\0c0Q3de3TL]B_HCc\0ba<b=PIGH8L
/B_][D<W?)SP=X@F;8@V0cIEa=)B\8/-N=J^:dF:DK@7QQL_&FGfE:@LcWbA(^RB
4&eUYR_S^>:AGF3eJg8+3:59CVJ-1\Ja>:VRd[YK+<7VBJDX64bf;_bL8?+I.&Wc
_b_25O3T,X09OX2^Q15KPL?P+H>2SY@,G7+IJLAdKBQ?C/S3aUb6A/&^fI6F-gR5
CY5<H@5O_P-;R;VG&\@I/QC<?+]?.(G/RT<Gf8a4KP5+^V.YMVA;6d4K:_L@,OO2
C;#>bOS)O06aXcJDFN^@c^<Qf+7;YJUXUG>6.P,#Z0aM8H2]8(b\Dd@39NV1=A<e
3-gP_8RUZ2_B7)9Z&87ZY5^9L8Y,O.6FY0RfRLb<JW6BY1Z+5CHP(I/8-e1&\^6R
@B#8.A.9L3V3\40D,:H,0=R(Z;e8@LF#K4gM0+)3.7FWXeC?O6gJ]X>H10/K=BV.
b<H[KV)0[M32]&,(;DFH1c#PO3/(DAaE\GD51\]R1(:5,\e;X)O?:NURRKMG(+U-
S>_-T0XY47=g1_[7;7D8GFGD^B<.L_U71\5<A[;P5[c=5SIFD89X6Se8RJ9H8Q8T
KA@JWP;L6;>V&a>\1X\L,bU-bg#EOHTL\33K<\B/+/0dMWPWe;1=^+1f8McE\-;c
HbM.BKM>U[RDF&-\Y,E(J8>UQfCK52\Nc.8b>X3+?@FI2G0]R-Y=S7W2C&.ISMRR
Q1@O+ED#9H:A;F2KO+BH7:ZgYg6#RSOS/@+cDA[L@2:bK5:ER:[UMGC#XF6Je@ID
J9(DLe9[C^=L=>0;>(X@X1-2KWSJ.+K=I_1BHPMTMUN?&<@<\FEV),+4FaFZ(aB&
)@4SI9&P&I&ZG)6PR:=+ZYKYe5_Q9^_3MA7Lg)7T^LMJV-9<O6P\5?XY2E4,;10?
45#L1R5,,<CKT)b-(S]S^eZ&>[d\ZOSVCOH6C-<A>b)-OA=^]KEJ3D<<,1H;?a9J
=G\GC)L/G.GX^3Z-bL#Aa/D1(c@>T4[CSS/1#IcV<]V>Y)0#MNR\,L,,5gXBWAa-
JKP9BC32I3A6\+=fUggV[VHO2[HGA64McK+-a8Y/G)Nb^<6fW4)T7_9gXZ?LM-:4
Zc>X]VNE5)J#/FX&PL.#--[FAgWI9ca.4KP\OEb[5FbEb=YC-2&MYN7I[-:b7[Y0
=FWZd/b(>E@6]BcK,,1^=-\c[/>HTWZZ0beYCT0UXU3P]V<:3G;B1Be>c[D+TCCc
BT,RL?\:4A]+-Cd#-Hf+LC;\3\)(D^;902O-]..MQPJ03TQOg?D3B.ceW&_?CE@c
R5Q2fE@Y_CWd6QS<;e)B)(+@ffeXVGJYFZ\b6?AJ[R.bQX;K:ZA#HMQdK@S2&/S1
6)2cI4PH]YGCD(MTRWD23]W6+CN;N1#8FFLC]>HDE=VB[-U)4:E[;8]DX4O4f671
D3GECECDf^db?):9N)AcfS8SG2dC2-:ISVg&M3?:L-+daX<Y619,.1APR=AbDN(D
,OZIEL0I6:25R@DWXUDG,E0,C88H7LgM3^;I&15<g5)JTBW[+5b#\e1bME<fI3QL
fD]MSZc5U^]U2/IX7NEINaX>QWYFNE=7-NY0R>RD8d(^>B-M^MP#8C^U635#;?1G
&bPA&Sg-BIKdK3<R]V<J@DA.A\T_VH<2PHMCH47e;F^\@G;B?K.F5L;YNdaFBUKe
W+3g>_<1(/5DfB6a4D^,P]8.XNW.+C;7>c6_J2I^SYLZI^5ZK-3<7@6@M0B3:,,.
f=94QY=eDMIK\D2>(Oe5X24(V^S&\Ndf4OLfcgHLE8A;g2(>6FeR/]0f\]P:ES[c
78N;B=Tg\-HSSLUC\(3C8KgE-+bZTb/UJg,8-;5b^GXNF?\LaCZX6WWNCI^.R+NL
SJ93)]J[Me^3GPg2:[cG;W5H4MPcP.72Hd6Q12:g04GNgG.^+U5<WG>eBP[W?:BY
ffZ/W)GR<2<dP(ALNRB/e01eL]2+TE<bM<>.:#9ZYLCY9Ta/fK&8YIHQ3;UTH>EV
Fbb[0=0#^)X9;c=D+910=cLQbER5(/TJc2XV8L3DM=e[2LA\=VaO:0c+.cJ7-G1,
R_(>OVc^5116WS)83#-6PY\d&2ee?)[=/9IOJO9Td_fJHYGX@,Jg1UGF<9ZEI7+8
U:/;@]b])C]#B3GK[<a.)R?b7DabX<0O8RD@^6+\4,f@=N<3GI^cAO2,0MFL(A9c
La/:/ZFXXQG5MJUg0-Vc5@D([g6baL+M+Fc0\,c.[3Wc:bJdZEb<PVd0ASfL83C.
0CJI#]AfQE17]H1QRY(\ER^3P(,=aYN[,#FE.;1-.ANWZN85&.^4D>F9&AL,4(c7
bM,dHVNPQHgV,7RaS)N<c0<-&c[WDPWU4OC6a]W4O@G6:AM+dYW:>dO,[.WcG^a6
S.>Y#eM8EB[&,6>F.a@a@f2JNfH.=2b>[J:>Y-[aQQKR08+A?U;QL04C5aJMD^V5
7Z2Dd0,Vg=a9GM03E^;@ZR,]c+Lf>g3JJW3fJ(Ve&EdeM?PT4E[L<I_EgEP4bE2<
5U:,g^FF3?+1F=G1PLD6^V+NRJ/=&_QV1_>;Ja&:JF&V3d_C@/-fP^;53T.R/)9K
8OU7S>RS9OX7^53QQCBB4@1>O=>e6RcL;]VV(K<IeF95QJdc#(=S,fM8Zc1P,HgD
FR4L\77Pa?;9M:fT6B=QcO=O<O]1MY[LbV:P5Mcf#5P+g6=#2a=2PZ2N,/IJZUf=
d.SCU&?)Gf\cP7BG?Ab:Og);/,9RYBP\^6ICC3f@.SBb)]9@:;-fNbZDZ9C9AI^;
E19P4AC_\&d@1&EO^efX=gfBAS@bTbE+dONTBcI80(&,^#NC;HeHP3(1dEIGIMd1
+bG6T@a?b75>9H8<S^X/ZTWZW/&L58+Q<J28:;&,gWe#]Y.^[g84I,I]1/4G/QC:
X?O:#SU[Ob44(&J/.CC16a4I72,3ad)ZN68U#\B-_1BM=daEIa?Za9gGJ):AM5Nf
5;@ZD_Bg-=R,2:[Q]_^10-TO3/(1.>=#\3<,@=JaX+4gf9T^Ege:L:X7SDZc7]/f
DN(HH5e8;G1./[6^9:WXS.d3e72S_KcDMVBB?D1F/F=TJ[gFQN1cQC7F+bKU.I[&
2bICN0SK2\fP(1&M_P>HV)I8A61O9.;CLd8IP[GV)b,+<6JU,+OaV3+DJ-88X,30
53Q4AgcH+bIe\S>10FS=N6WEXOG],d4?_=8DPN@&@5a>fX-)#>aOe8^)OVDXS535
8\O3WI+/1JYg5S0-GAa\TR7X7RH+9Q?OTgPLb?71U))[/.Z6#ND^QES2fKa/QfHL
?A4P_/D/5APbOV+gg)Rd5GVZ3^(JAfH;GJ8(L^5Td.Gb)C/2&V:/9_^JX^HJ-gX.
^/Vg8+,T+<Z@?,a_X&S;X\8:7;-b/>J:WTL?XUA1&@G.DR=XTV-E+]O)MbUP0MG3
Xg:368DbLbC9=V(dFLbQ,/&+7#O7X(->&2A0dIQe+O;Y]>Y.#)RP=#@baP@E4Qfb
g5]<aI_O>(=_LTSSJ/T;ag#b#eeO,ACgPe?cWWTV-cO(#&;a985S>Jf^[1@H/aP7
aJ)_G2:9):fJTB^e#(-9R@))VYdRM4bQ53cb+>M#bg3R9d0g(N=2+AQNN22@2WfF
UV9b)B4A<FV6F],UGM7+W<g\dg&c39=OG@^QNg\?DZcJ[3[f,PP8Z52TC#HVZ;&a
<?-+P08HbFa[?(K&c6]BPOg_5PR6F>&?7g+6>d_?8P<4b<eT2X6\+AF7)(GSOS]5
J9fXJ7Ng?K?/H4RAK_MfdgB05<3eBU>1>92#URA+CP@TSUGCD;PO)\@G;^Q17-TD
/Z9\+Cae3\?=5>^)=/08,,H(Q,8=PJJAa&Q?]6f<T_/GF?Q&McCH\C/RTBVS#/C7
1T(B=R_>IdSdX8NL/A/R]9<B&A@MZ:M<7:0,VGQ\\eO5;X#=ZSVE9)>]W0[8aD:?
KEc+-UYK4W:I9@fe[FI[-R_e=IL].G.>A9g6]R_X[0g<c@WSL]SC+K)FM=<RX,F9
F4Va9/FCNN&OJg[>#8/4f_)9UH;bd4a[K7bHa2NDW(&8H^GG7LP0\;8YY]6YgY-B
?-.O,1GYI=67/VRg:.8&.<L&P_<])ZRBadZ6(3SG\K?.QUY5,5>X??^0NYWa0/BX
=0bU1SW6OFXW(JOI\/<M8+b@e@K([H)FYYNR_D\:EEZE-;5d=;/HS+1(L_]Z-1D.
7KIgCZ81#Y:XV81g0-[(FN]9H@<P3?a#0GH0;bca[7f.:G>TB<[dREXG.[E_Tg>M
>I97#8V#<b,E=2a.ED0SB:.<=Ta[WKR-I7Y29)_W5.+#R7@1RJa_R6(5874Bf5O_
+#GND>J+DU)F)2#TdHYdI^/W]/0Be2B8Be?XVc<(96<XZ\ZCdTOKK11SPS>JO6:e
f@&JX_X8,R5,WP8+D&-7g=G52[3Z,1&b)C3M7BAe,RZ+XY7;5-@/K[N:,BX<8MLZ
.S.4INU[>BO7ed^\T0>AN[/+2=0TO,[(63]VQ0<e9BV>7_J44HG^OJJL,_\R:ZJS
f#QJ54a)S,cT,F4\^gD=a9D0N-U>;^?.5\RAI<J@Q/75g9GPPf,3Ube+9b\^KOgX
UU&ZW75^EKA75-Xg(;f31>CXZFG9UE<.X3ZK-#VQ_8fA;P?:?eU:?c9(Q^IA7MJ4
<L#T/^G536S___(JL:0Q(BQXgZgeVabPP>81^3B7-\39Fd22(HdDPE=ZRD9WDZ).
(4O?aDOOCNX9.8U1dP0?FNRK\F@W97N3MDAa3KY)f\Pb_EEd)W+BO77^D9+(e9=#
O&cbR@Z)B5VS4AQJ@YXYg1B9,49g64CR.,ZYO?HPVWAT)KK2aMJc^:12@&+6648Y
K&LVH^aK&(JLRNZ]7bU+X_]M6G]M93,7(-;b#;8gYL,FVF/.JLN4IL2CV83TGT.Q
:fX1];WFM7,/ASG-_^GHXSC7W(7H9GdT>YG-9Z<PccS@WEeX-YV.M/58GK6OJ?XN
XWR:TQFEME+<aO_3HGcW>Sd3M5+D>,UZddMNYT--O./@<W[fgMa6&Y:+-?Zb<0J^
Yb&WdEf5&QH)GZNa[)MPDJGQ?7,,4-7B4@QQJXEA(#2e47d[b)[Cg;L)PGTOQA1:
B.E9=#cMEI([&)5YDK3bNOZEYZ<ZD0,XNC+2C>M8Y>JRQH6cg0a1K-.Ca<LH^/-H
WTfTd;=C33dZH_WbZgJQ&I5SCON>dYR]KQKe_8OfNQA9LQ3GG^41]cY<SF(He9Sf
07-+b5.J/QIOPcE.OFUQ\D+UGQZ5TU_3BQ=U279SMAfY7^4\2;Y?[I?HM,X;#7[Q
8&_MCE)DLb?#Q-a7R#CKZ,L]/fI,@/Se\S<PcW8X80.EI&eR6&AW7F0FJPRHO@P4
2X^EIOgEGT1/5R&@J;9O9#:b0W))e#/C>2+-[g)dAZT]\D_F<MVDQXW,e]YTV+eC
5\;P<@W>bO-bXINOHTG:(6[JMLU;7:K2BLX>CM(7S<c.Z9UT)F@Y4JQ>BH9R&=dU
4g4XSD&J/\RN0e1E(Q,Tf6HM\,-aX?KfY41;&[K>=>V_<;21L+09TNSOH)_:,-5R
/&5c-_J81\7X/8G,OD0CE>/;_\f>d\5<;SJ2V2QB=6FOTB5:1-HM[S,&2><T5Z;:
a)gQO>.X0Z?EPcfXM8Og5&EV0,ac^N:OZ9f))a]2<,=SD?UKD&bKg@XX,b,&0I\>
Ee9OH-E.;e6(MW+(FU89QCX)JP.fDP<f.J>4]:dcPRYYWf5b/&S,HT:g3B;GEK6A
G/aWFI8I25-<@aMe_RWaHfBZ_<+.BRgP/Q?LJbKY&=.3N7-)07@,76TIH?KG&>bb
G&5HT]UWg&1e_2F&431-BO.Kef>DWfOS7J0=eE#VXN9L;fJ]NM=K2a<&V@YP9@_:
-&eR[bZ<B)a?H>H1fUB5-?#]gAB2E7/aLP1[H8KMDZ]T5F5eISIA22g^JI3LQ#dF
d&QA-Ee=E7=\<\e@-62Q^Q4]D.bYbM<_/dN=d<,KPS@GO#5TDV6Wg&Z3=c3MK)]O
4H;PHJ/Xg]@_EK[SONGZ]c4dN-C]cY3[<X91KDOdTT]H8.#N24ccW?La92U86))^
4_#8LHH:fPJVa(a^90bGL=Y:QZgZMO/?)UFD50R\00QA#VMELN=E.OEU(SNM=9TA
SJ.2>NRH6RG4a^f-BXe3^G:Jf65c[d25H?.@#TOf\Y@,B0[&G,3-g44WNRSRg?IL
3W>8I^7bA?(CEQA7&;a[TC<dPN4-g#?UCPCbFPUB]K-)b-TU-I:d]3e;)A_6H02b
_NU,HJR#GVBH#CI>#]Mg<D-[<bccK/8MY@Z0IO?P&&::^Q/FLA.+Jb[g)F1.bGg2
Zd26+6fC#IU,155,^=6TY@-5WI-\9M:Y-8>\SSb7CRJ[.g[9gBJgG#)9,C.Fd1D3
3FYC(=QU8I;:14F5Ee-:=eKH3ee5M[WV[]=:VfH1Ig9Sb)V9O]eg/0gR<@Ug#6YC
.-0S>-NQN-75:@77QUF@GF[,5WM3_gG3fg628-L/)=Z/QS33HS+=_[)gUIH23_@B
L1E?F7]R5-==+cRO3=aD?dZ;.U&>6_dD1\65W4fACEXG7NcN3Nb)2_Q]?K0)0FfH
[UaU>D3:EB+N#-)5Z_.F_SVf--3]D.>Z,C:^DJdL.0[8Q9OC4YO,::RB5=0/M0;1
CMH#Xd-4B9RcRON31)3MS5:<P[?3U]V+)Ua(1GV(4:YK>RMZ/#EF,>UY+YeL,-7Y
<Y3IG;0N8NF7P<0Se+b?ZT0/YXN6;-U,TP4XHAH4SBZ)f]3<A(\)L<:2SS0WB)=1
@(-F9PUW.KfW>2>2<Q53.1MAMQURI;IJQBH7S?+@GW^cOAH+d8LTX7e[a-()@GP-
e<FN(<KF46cc(_FJ0Na/S+0bL;?dTa4dW8(/Y3DLE#/_>[8V0Kb(XGV&D<=8X;S5
K).+]d2OS93..DSf/U)g<@g?BVG^dROQU44F4-b7Y)fMfKV@G-5FVTN_[SAMTda#
5VH15f[SVR)I?>X5MbY[=PR^Tg7)#<6ZJ&C8[JbV6/X(5=GSPab^F(BPCB[5?N\;
2DaX>+0:G]S3gU6?DgS7I_X>,X@f+dXEN.AV]5GC\K^e,-[CP1];:>g2QZcK7MT4
cVB0=I]9G).EOJeC\DD?7>;&c\.BO5N)2fF/7+Uce@<2/;/,0cbO@U@U].aQ9E-X
Lc_=01=;3&1U/FO<_?CBC:F7KYgX[IRZRZL>Z+QbR:Y:&gCPBNMH7SH6gZ_gV\IA
C?DD29A);5T3?N#(JSFZ\Me2.L>\K,MFbXP#5M2-UOMW^;N[DG)W5/dY=5^(/DW.
a6S_=e-dAJJ4f8^NT,@ENKPI3;.;HA;)01f<I3<J)b@DL>8+&?9ZN/-@#XLc#H@.
IEQCJBb3<H(MB?2W6bF&cc?ARC&S(cD<8Rg>AGWU_5X,McD[:6Z2#2_^,-M3N<[F
aZ?-SO0Y_X+aHBc=0P,L/O;H:(OTL-^<3-d<8Xf?[EO,Yd4VG=OOWVUVKbXeLIGW
HG@8K0U:7#.OH1,N>[Bc-[-QaXfOEZG[C=@\5DGa<b(K>9KFNKQGVL@VU6[9-OON
VN2TaXA+]3\8=P;>G30HL?;T<<V]?&M-9+>4KHW#B@_07;>dDd+e)X=/1]GLNb)@
8/QOZ]=gM1.RO2.26EY4BB,&H-KDgTb]^#+6CcbSN2HOJFa<>0P3NTL/.e@-1)d.
\KO;VYEG>:d?<NN>,Y9KZ,X)KHG>aSX7&NCf]-V:Ee#Uc@;Sc+,-Z_;7AS&E562T
=@_AUcQIa_F(]_)>NSU@L;P(MT;Cd@Ha\E(I;W7.UI&fDY+2D_7:U.,e.K6G5SO]
2gPOW6QgfdJPW&&:U)BA,MeXK;?KX7;:\3)0F9AV9KWA=<D,<E80ReT[(b1.;TCL
MJDON.UH##\/22E1d>6fQF_Z.>,1X=;BB]VEXIfa48f/V]V4;W6#\f8aDJT1.af1
,V2S2A-\,[dfD9#GL>BJ&4c^0328?0P6S:3=[3,S@#C7S+S5JU[2c,A0<F3Q5Nc+
U2VHWH_fC8X/.1BB^P9>;).c\K=:PYTCJYQb1#/9M+#GPF9?S))[U^;S;\9JNc]K
+<ZUL@=H_M:#7FWXE)4(,<7]b0:#JW6HbU6LB^E&:D/]@3N,d4_FFdNNP=\)Gc<O
[_<9UDF)T#25eD/S^/]TN,5]8:F^5#gJZ3]7^2LWC0J(YE<O:AWLa(Q1Uc<W^.Q_
W5^)/A=I2#>7Z(SL2?KE62dG5L;.Kgb@X3M&6NRLI^^-_/4e-@AIU,dF<;f0LPdf
e(H3>9]F8JQRbOX:8SP>=ZB\.A)MZ#3c.3b^NYT;#3eEJ]@>NQF:a@I<TTZfLc+e
=0bY0&EVMf7^GF<b6OXT3<X309@2Y=I+4;QO0P4=QW^<6Ve?58fNVG6Q@_g:C2Ca
T;g-_@_/HY2KS_,F0Q@J683fUI)?.G@KgfJ+LNOG?];G.UA31Ng@=CW/L0M.,(RL
e#gg#J&.]^N<44JKb<=G+.+79&db4(Q)Q(+EBFd8?_B3[NW9<ANVcYCf25@80CD4
T+_7:,KcZU+6/T&S:F?c7-f#OE7C,V1-9(gW1)<A>+=WFdT2MLN/8,Xf4+<NU?K0
2M?N#aC-8\SAVcE41SMYB]DX7/1-_N^+RU?GT7Tf/EP_G11>)YJQYG(63U2O\>6f
TWc,ML-G[1_;5V,]dK?Od2WVJR6gE/^+9L0)3XQ;a/++cOJ-IT[BXgA46<+@TP^2
_IV@_JQ=D3)d@9\UbMG1F-YG&CCcIH2;HD3FAN2[9^EB[F(031(f(e?B4[KG=?aU
UAZ.WI6J]1gJFfXZEAb2YV8X&@C=W(GDC6e99MELKJ>P>\J=]Y4D0&Ma48,D+HNL
INFa\U]fA;5cK]9a>)?Ng.3=/?T;@2K<0/638.Z?5[>KV_XZH9eSa4fD1XO_Q(^<
f6g^[8NN^d9WQ(K/\>C.;0-aGA,3MYK/BcLaK@7HS@F5.&b/6O,LUO+XE612R25A
c#g;<\cF2GILHA;X4S-7H0]9R0f.CRI:V]I&RT^WcVQK7S[+WgaSX8(cV)IA8]-P
e:M(W=J1L&W^A>F-79#X7F&g#SSA>SP=a4CW;OdeS15eZ(=KbFPPI[ZT@Z3\Za25
V@-[2)34_D)gY6-O+/2024Y@)@:95Ef)O<\SIRU,0NT/5:cA9IC>dK;dZ\KSV2+I
e3S>d^3EJIXC:HbACD_46VI3UD,67@LNM/<JV00:V4;@QM5N>6H_d9LY<#8\PAC9
I2K:PPH5?CNRU6bK@I=_UdUXKDXQGM<[KQ?7e;YW9PM@>J0Q.H,^9[3@C(cK5TT4
Nb=V_Y-SHD<(XcIOGL:Z+bKOe6P#R,4;)O3YP_&.gJeYc9PHLP5?2X1&#E<Q-K87
E&A?KI[ZI>8^_4]eF&K=9d:Q&SVT2C.g-2D7fU>VNBJF)DDHdfBa-CE+Nb5<E=W2
P1HN+2fA[1\CR&d\5([&@LbHSE6(,Nc;U[3RcKF?ed5YMKFBADe=J)=GP[#6AU77
[7PISd5W9HF=Z&N9^JN\6_;]NKU,]&CGESd2\<R6.[MYDX[+Z<Q1#RS=U,76GX4#
9@g[@ccg\O7fLLT_]_e2ESaf?HEcG5.B4JYQE+L@3\Ye^70eX>-18SF_b\(BUJFK
;d&_IB^+1@@YBQVGMK99@-RO,I[eFe(7S&D:@I=W8Y]R7(0P7gFe9_K_<GA/VS.1
(DV^DJ9?N]eP,a]5d\_P=R0@V9(S(c@F9fU@H:a/ab(X<Z>R7aGdHgdF3F[&Y5L4
:^ASIK3J7M\9[5DR2G=)?8-DB20WY_c_\bPS@2YJ3\A?LO)>+fZTB&USGM]Dd@0O
[U:WY0bS3M=Y0ERfICJbWJ_BMGPRL:9,C_/N/]260]fd=GTZVSI,OW87a7TI1&H^
eC/UN(7?g(C=FY5N<G2WeZON54Q8&HdM]9)_6_</V9:\b>^)6F[O7Kg\eIH4g_3/
V>X^2ff>_[OVFR;g_AZ+&5T/L/^&^RCP9B>a)Ba8d+BSY9Q><ZML@#G0MS.fD321
;f//TILJ=:UH46=dTW9GLN?GZ3LM,b8JLU,3#^^=P1M(U2SaN8Gb6HM1SK7g)]WR
S8:7//RX:/9SJS\,O9M&#V>FRP0PdafBbUCKZ<0^fI]/KZN16NBJQ+_QOP^,&[8L
ME]KH_-6PdX/L#Ad<C2a8Q3fgR8Y53WU8&Y3F]ARO<LS2-D<XO2=fgdK&5B/bZC7
WSf6.<J&<Z_.5/e68O<.4S/#&PLebDM&H+[4DCFOcWM/g+Na2KA>Y?VP];NV@6,>
.7.<[SC8>NW@@?b7J,S-@>f&(b<9LJEXSf,cG9+F-AZJISaDf5AaD@d07DL(=eU3
R<3\3dD)]7Q>BN_]3?JQB2]a1,55IPC,cRC-RK1N9VPVK>[gV3Ff0#b,4//6:?L0
1S@4-;:RVaC5K8#fc379A+9J:EQ#+76)E#e-/bC36)YO]79U9R7Wg.N[d.EUK^O]
\a2;b.a8@MTU@@(/80_,@dKQ\1dVZ[N]aL8ZD)PgSSE^P>2RBeDIF,L-M7JK20Z\
##BEe]4Q85<[=3+SKJ-56P378^L;_OL59N,,DIXV8,X+;^CgS[3=HC&7GQ,LP0UI
.JafFBC_J0VC0>B_84#=3@2(^:RcPNU(D[2gEc&4I9=/bOT:#H:KYMX1B)W7AO#M
Yf2ag7^&.0)(A(]@T<,+568FYG-+fdL;C8/5]H6\Tf_HQ_Q7[+IT+#SSDA0fTLJb
33R/SbTHd).aRW];-EXW8I^/SV_C@1+NTZV4\??E#R6deSF@_gJ6>W2\)c&E@3aY
FHLFNQ==7,L\d(Ib&O^.[E_^1<G+Z.JQPYUSBQgYWGMM4dc)Hd+G@DMISLL,0P]R
T/TPV,@2B49<Oc#[KgPK:N?CLd33:BJ<T#QVL8cD\Hg<X+g@DDBBNDKFRT@WGQ_8
+-N,;E]P&^MLf+Z=CMeeO<38>+@6DM(Qf9QZKb2eC?QGaS5C4ZWd5:>A-?=@G_/6
P.<efbGR151OTG4GBK]T_BRf5)@.[_b3WMNY8ReSGT:Y+=7@MRTC-HQc(]]F5_T@
S:)8\9L\,7NLHM+@d#:9SEf)MAGWY1A9([2EI\@WAFH6_H3\+ACc,ZJ&UKVX3<T7
b53,,C&R#L.E]NCTfBGBB1D:EYU.PX.O=[\B(cRbaN^VYT7[E@H)XZf>Ad?)e:;/
0B<[VI#G6UVYL8N6O+<\)W1E=&_?Z#VDZEJ.S@ADWSKZ<U6S\EZ,Zb>;^2^Zb.,#
[B3fGcW6c.YKe,]F(:.BSP=N:RAN)XI?+Y9W#.847Q+;TVe//6X9#_T:T#ML2=/(
&2Z32eJ7EB+LbYe2+BdJH?C3G?-0;4,VTXY)K<BT1Q@X:?gZ9.[[<HYH&</KMF0H
RNA//J?a<f8DAd+PK2c1c]\2@;)I#<5)@+(8DZU^FMIM0C)5EIaL_[)UI_:VSYN^
L\^T/NJR?^C,gGPY<UEXNSTWK,M^487_.YgO#edV9<\)Q1-,O40IbQAaP05fCTaS
_ITLYdd_bb^HWRVTf#TQ2YQH5S3aNYU).aB8=;;R35,<Z9DS)..Z<P1MfK24VSK,
-aW3502IS^B4dB^9WYVHSYSb+?-bEMDQ<E.BDW#6;6EDGU+UDL8e6c^?H5RBSDT=
=K=Z?+8NQNR3@9e2V=_C5HBN/T2?3/GMLdXUD_H740X[_TVDT&>BEZ6@084CdO60
+CgcZ]M\Q.5CWXg[1+PCWaE<W,<N^<-4@5&WFO39/VBP\LLG://>f3^U/f@#YXKY
c^(UDY;Y?C?Q4179b;B(Z]a//6.#I9feD;PREE]\^7\6,HRc\5cDaXS^37S_T6H:
FN.8eUD1[IU1XS7b<+8.>J_a,:+_3(/gf)1QRO/FJ6P8:O.(gO0Gd]^G\LWTXd#Y
:A&.7\b(g#e2PbMb[T^bALfda&DC,6U=4_/RAIM6]gR9eFAEV&E_YG^U&MP#@ce=
@L[Rc31O\aO3<,3ZZ^U:U^S:2?9[6)=+>Z0/D8HUU[4?Wa#0O^;L^BdJ0N9>^K3f
^O?B7W>EOU[JUf])95:7TO@aYgf(8[I>SbN1<S@@5ddcA<8D5K0>^GZY.bE&MeIT
)bI;;b\S&5]6).VPW,2.YGSFSfK9J/==0\J<#I\8)^/d\(:_bOS-PA70:[A^Z-Ye
T#YAd(TMLD09<f0;(H<[[)J^NG=#KTVFMXbV;U]Hd&=+B>HXc\=_g::eBR=2^K,V
fa;ZfI93\X/CC2ZBT8=;Q??F7a0J:KJ#ATXUd+S]NOf-/b[FaO/a1abL1PgM<].B
>&5:;D@2b_9M:J\,L><82e>[I<(HAbQM7/RefaGQ>5AH?L7<96a=5T<N,R__JPQg
Ie&bAZZ;B&5@bJ2?S@Q[@Ue;bO,HJ27Ngg]dG5c@XJ+I2gM4SJN_](<0,U=F@NGH
2f2@E0a>F5?&c?c@I;C]R=M3CbHDMM2W=CCA1Af7;#HUD:I9.H]Z84=E#HTdBgP.
?SfNBO(O4/8_;8Xd9QVA,=#^YY0G)FFL;>P;_(C.f@g96OV:ge0RFA,;+#+WK(.\
:@<TcCEXE-4MEQLgPG+8Cc/<AF(S)ARQ1?.c3SFP_a7N+\b2[&Q<CF)>/d/O1VU@
5:dD_a?Fg85+M9UM3TAMEX@3^29.P23bS,NH#LaSHb=<B5Yg0,P.aaV@5JaEKOC?
A2c.O&dI->;#41T(#<Ef_9FV3H,3Q+M1=_DbbR#fOA/)?GR#&CaT378gQg(a[.#K
?_XL]NOdT/LT_N#^?U2,DaT&>10WP\0QG3,MC4P#2J2\9<]T;J=:D#;=4E2,?/U=
/#TGD@^>AG&C=8HB/OM(<H0.aGNGBgTY):.FdE5<(OgS2TZM;G;b;Z^07S@fCe(Q
OG#EF,H/9I>_FJFV-QW.H2L38N^/gC-T^YY\G]>7GgZd]7f-YHK#fQe#K^7\W3gE
d/R#2@@C9a;H)X_.NXBGDgbTCNP8U&WUC>gdJVVWBA&Q41LaJ18P3:G2Z.7g<UX8
/8L&O[F@3#JGZ5Z:YAW1WR#9@P=Ld^cM5=d#c^9VK>W80GbW&;8FA2VS^:QKWaB1
AT-?OL6MJ47S&@>HeF[H_2M17baR8A4A3A9D2Vafg;3-1&L>OZYfRa1YcX2#X/?a
:C)0LO97/TS7/J.^@H)ERNETd/-FAE6d]TfMI6+3:73=f-4e;Sb8D.(JgAS6dV:,
?fOEU;GdETS?]J;^b)1A2551P9;W#DH[fXNJ[OSGfP0+.&X4KNK[O&6Q_e_2BNbY
fZ5GE]>V_FMaad)CAZfU6]1;XPUJ92M/DFe0S<UJW@XAT8[=d>3ZXC\PW8g-^,]a
?dbK\0X\[>04c]#+>/f)bMAAG6_V(YN[2G<JV4PJA:b:Wa>1\0\DKD(UXVBIX.[8
1a_B0^\7ObPgJ)ZDJ??PD?<Nab-Y5.a)7WILE<66f(8-GBMM4E;8\R83VKHJgZY]
7MXXHdFYQ;1&c6\KU#K9)^R+XF)X7@APDT0A0KO;_X6VT2P[2AUJfXG6MZXT/BA^
^=66CGJ)3D?P)#b18dadH-Q9g=-_TNe(XVZCRc1,(FKGWCF7gfR7PRM#5FQ3Ne.C
=A2NJ-]2AP^?cT..J^Pg3^&\Tc665H95AYd1EW9IY<A?;f034BS.CNW/8:6M56;/
LKbOAc51b7MY0F\GB3+6UX6G<A8[fQD_14ARW<::a+;Rgf9/4/^J\/Y9<.Pe?#-N
=62M>-dS;eIKb9R3:B2d-.cGU+gc2/HP6Q=7a@Uf]:Q,9)f[JUb)@+LI3aJ.K]]G
b&60X93ZWYZ+-D&GNP,cCD8=?_Qe<U/8HGY_>9A(+dIEWRC3b=[[)fd:4c[P7g0a
MWb13O/S.f&JK8Vb=OQE^IBTUBS=(?;3KCg.//T-&^NT-2\ZMaZV\/5T\XA;-?I5
>^0[F11AI#S_]_ZA=Rd[b@Q4]G25fedC5\04f<>\A5<[FSeX6CAL\e;cMBL/c)+M
CO3^9.2/[Qa0DRFIVJ=Z4-;\[9Y;JbBBEP3,\#_^b&XN-K=D0&P\M;M>dZWK7^dH
c2.\CcKeb#[87eMD+AKLFS\HP2GD@S=3UWF?1[=AEI^TCDS60e?@&9Q?_.R-G8bb
YJ@[(+R0[0.-Q,I5:8@=^[5Z:P=AM\L/9417f2b4_120GX3=cK_MWAJMWN?QL7/4
(WE.37TB;H5C;77Q#ZSF3VMfa>3;SP(Qc[(c8cV1@[a5c0:KY9@?Z(\3c3VR=(eF
O+3gGTdG#[:&4ODEH?Z)XT\#aPC&fRI_>I4cfF3;@?68C7=+fOZe7ER:?U;BKF]6
KX(JU1WI##JeF43E]KKg44A5(@e^52,]O4KeN^]J6@_2G>\=/[E6eG:X.,L5Z5VP
c7;IL6V/bMgW+Rg(9C=4dUVWHX\\=NgSGWW3RPQ//1f),Z^Ag][AQUAf6)a7ANc6
f@Qa@fLd&eW-U+RcM5<\0VMbG&^Fe@BI-R=9E&C[2A4)-PV8cd;fXT12A#\&cWJV
_8_I57(f<]a1?6F390bVR^6?4)K[J?BLJ=X[N,dB&(gL]^DQD#LYXHP;.?C)8SEF
[Q,[FF[IPNI>U:MRY9a<3<D/Xc0P_WM58BD&2;CE)BV#]R20;#_;4a=8K1>JKLV^
+f85#BYeN@Q:?H=HbTR^\F]<R6\_OMO)IKOfT5VT3=LV.b1X[8,Q,.4cU(4=Xb)(
ALE^b3:LFbD61bGHA0aN2eGIRc/9.D)+b-XNDBZHRBVHYQK:]?^A0[O9\#\)5e#4
V&EK;MdeaOb]/>S8WXQ8,USJC9fFH,gT=4ZC9\PW;B6RRV1UC_V,3d]Q2JR(Q+JT
[Q&0#JHU#\><T(0SEa&_.)42ZML\CgQ:gMdZ=_dXID+TL]\R=;QY95[B_b?WA7(&
MX+0,#d)5P789cW2bc]GeV^7=K2\BZC995B0\MYX70GY,.]_W,&)/TdLa<^D0VcC
,WU]bEWQd#)6^2];N;Y<YVRAY?>((Z5PXed,+SFP/MLYb1/@a/PE1S48D<;1(.N=
G)eM+K6]+@Y-MXJ@1BO#,L8K/&UJ==C0Ub]P2&R9XU94I^WX0##ZKI6R,\FYM7NU
CHM4.B7WN-3LD6e(ObVAYZ<1(O0\.D/@QK1=c[dX0&)-WK8:>?4_PO03fJY>K_>N
B@KCV]28_a>N?N9^J=DYf\IK<4ZY\<_-GXY>DZ^9gO?IMVT(LYV-OOC_S@&<Z0G5
/DR&_(VRAXYSEd.M])BI(D<S(cGXcgDOXK2P3IW.QGE&+c0aCF1cA2ZP-#c;8&>;
B;K/_.\-^KE2BgHF-?0#XYTWWBQOV#0WY):[A?E<)b)2E3JD6=P9I>;aA-J?0X(2
UA>9acSWUXSK_A(K15AUGMC.Y>Q_J+DTfWC]b:K9fB^CFF,L6_;bTMfZbE)G2U??
Y\I^&OU6=H>P+WRXMBW=F;/29OI=<TcF?P#39/OG?P(MF>M3H(L:WJf.:\(AF5Hc
4#DK\Dde/KBdef^+C3+NI;[+=0^[O31Sd0.MQ_)JL:LL^e(fFR6Y\[H,OB&U1UU/
;4#MTHX^[PV-4c^fUSg4M3)/UIVa+Kg8B=Z7-JV/6Oe4KcJ0Z.<L?_Oe5:>Q(OY9
C2(D:SJ;_7AU1Oa/TC0;I36[)2O1=MdMH/8\/+g&OFd_35SR2CY20HgM[C?UV384
5QeY+WY6YN]MT_DK0>@YA@YY:,E.Z5L)b,U_XNTD49M2ARfYSgUY\XF_aM,R9WY>
U;S+T,,&DP15K86c/::IDYS=RgR\]\YW@d-d/4Sb82<8gP#CQ-,T#Nf.D0X^T@]4
<F0EA(Ug0F\[W^cc2Sc)EA1I_V28F3XUN;\]_[GGWe;PXK.XEKB)e>D@dGJf]^#&
,^L20fZ;g(3:3H0_7VX_Tb^[MTC7Q6<=FNFg=e>K@#S\aQ]/.^0D_d(HP?Fe=;XR
7T:M8B6+Zd_O#27PV?;_S#+XME3^S&ge[3A7.U4,L3>O2T?5<;]84@KGb.Q=#-@G
R0fZRK6X6E/:=OAW\@6T)&cfNJcIB?U)[6?=R:=_5GBO._N,E)KN1[]VF@;D8a@/
FJQV(ESb39R\cRIQ1&<3OAKP=_6FBW[gRG5A=OdLB8eI8U2d<LU9L,_fN&Q[eZ[0
(,UY<_8WHHJOKKZT.416MP8(O./P19OE7U?=YE9_SEBL=TgW:SBLQ]/SSd6Y&0ZU
8Q7-+b<#AWXS<[[(?DNgLJJ@O,.^/(fFJ^WO(2V([]ZLD/.;#2Y1c=>79E<2T_;V
EM7P#6H(&S;KMK-9OQ&LMd#@Q\Y7?HcU3.\:E3/N^,5J#g@d;e2b9=N@MA0.[\e3
Z&Y6d#]JRe,V^+Y8)K<A)+0W5;RQ:R-?Da+8YEYQHMNLKWIXJD6^CQC8@Z[fS8ge
N]54M1Fff=EVU<PC/6F<(g,<b@Q#:L7.D<^D:I/f[N=](-e,a8Z+f(:c(.,WI</P
&+YTM_&\aaIeQKO^B8?K(\,XS.^J.U](Y8ASf]=dZT;RNbQKMJ5<FBR]CUK\-a6G
)0^/(^7TeWGEQNXOS5g?^9APP5IG57C4f6L6e]F_aPL)0f(C0^;NFB1&b+4?2X^-
I+g&9]=ZF4CM[UdS8^RUC.G:&9,c^I(7T6ST4S/WU<4Q?E9JD_0]VSK]&PSNY?RY
M&56F;<R-Ib<TZcXEZ=QC0+=2GF](YE/7c6@dX7bUAUPL^FdZ?[MS&<M]XG6W;BB
N=D:N-a(,1U[2RaU5.\G[T.0EVEG0J>J?26Z>aB<aD(L(A-\TFH]3<EBWUB?CR^G
84=Kb&XKFABg+^^f=c1bgQ@XRB:]&dZZVE0B7&;MV<KFQKHPbJF-XLM2,g+_U-U@
7SXQ^eJDdK#=-CV:;N14N1(f;]5#N[,-<TE)F\67)].DO04@Se9CKSMg#G)TFf7<
\,0=)QC:d6Ga0-M?aaK:E1+f7^:H.gDX-fYM,R2U8aC@eJN_feP>CC^;9X8&(8?S
d;?3(6gf^M5eCV:4F]67FZ)cCY.K8[51)NO>aC5dG7#]8+d()<](-eSF#&;YF9MA
QI=4d-2Jg.-OgVe-K@DAfN/_ZD[I.O;DQD11d^?T9.[CRE=aB\8]g?SS..(,UW)d
?\S?HQc73;9/-9KQ&@6)eNB+d)E?_GV/;I1^,:32VMF?cFQX4YXf0KR]\1BHVS6Z
FXW,)abb+7L4?1bf;8E0#S[^4PS#E2::XBMf<bSMcRIe9Fe0N1MGSXK8;W?,O+E2
:Q5#FOR4aP[169fCP@3S)#_dFg^^OYS=B8D1\JCB&f12I>e^M])2ZO\+/<0bcJZ5
OZTb>.IHa)HBY+NVAM4[gf2J]e;U(++M>3?<6)</SdPW,:X[?-E,R9VY^eXXM)E[
PZ9(f27?g?2\]1]P&8,\Z\T1A#>LdK2BB=S=Z]2=R4@CXNGP/][GbcaFa[O75D6#
DQR.F)-HBJ>[^;M[^=(1J]ATV,6deHeX(CB3N86cV:EC)X<<F#K?6GZ]RRg9,JK[
Y\.R:eXDM^F(];XZXV>K<cJa9d9G+HXW#(g1ND6U<aM3:4e<>0#Ge=IgRa868_(Z
PU2MK_L5b\N7.7NdF[##0Zd2_:ZSC,HPKBAa7Z(0;@]b;HB6BS_16Gf92USO65:E
W4LT2a3d\L\(LB)U)XL3,X^0/Fd6=W_@dO,FcS5JfP#2#JBHUYE38.1?1(R9VfZ3
EFY_TA9J<H.PZf-=A;Lf<;:7\M,QQa8BVR,a:0YF>/d-XLH><MF3.D]G.NbJQ6Bf
Og;b:d?2Zb:/[b/R^gX1+S1&JdKJNTT_Z3>Z7YO7_RYCZ[-20?HGcQ>VYZ[<+-.:
N:59^I2K_4aOa(LEI+DN&I:GKYAH]TPb[:ca,Ad>Kf7R;+Ec6]RK[_K5C=JScg1>
>eQb@3W,&[b8;O(XOLaF_:?WdIJ7<)DK>EP^/<1&aZ<VDA?6>\S[A1?2I3,I90VX
M3X<JVLg8>,N4,9[LH=\QPLL2RQLA-6TH;Egae,c#RCccK^\8\+(52G-gN]B@C<9
#1.b<\dc5>+fS?GYeR_=26S&7#L2>D54/cQZc5&,00U[X49;)A.=c723Ca6.b<56
_2aB_N6IFeNLL3L8?8\L.3]bCaVA>SAC1H@L4d2(aX]Fe-UFK/TVQ31_a]F-d2&,
6(eNFCNUNCS31_X>;5.fYMS[1-]RaZEgC6N+J1#F<4=;Cd:9JB#P&^97MT>=#\8)
;##U.UcA\XQY[T2:8cEGdM1A/cHB69&V@gFD]G4K>K0c?=G]-7A8/#;]XF&;_b[;
\[EA0CN93H\?I7]EY3>IZA:G=3L,CZ25U=&&7U<[b^(LJTXV/FN(0KF>M5)1b[(=
H221+]4F0QH>g&,-fa4[&+,gLf#8N5\S2H09dQXaAb9MU8S5GV/QWCDI[-KEDYKE
2a[?814UM&]XR0Q.E@BYbW-Y,AX\_DOB;F0X9TA\7cT/Q[DK8bB&<1?A4_(1]>2J
cQZ8,,LXUJ6U=,+9g1MP@>@a_^&cUCT._K[F>Za/LGeB3WGD-U_V.VeV;c3<XPeL
2P1UXQ)CdJ>\,94YdPMZgUbJ?YH/B@MF)[R]>4;G?YKP?DTH\+4<?DXE@BV5UgKA
&J1H&aS^9JX/b>F^6)TR6LP5Z&c00Q572+Q_A,&AG;c45^afGU_K_dN/eF-?gTA3
a.=F&<?[KYZSO8ZROZNUa8L3]4Z:\&GC5NH4K\#,O8aBFI0\+TL\AC2Y-;LDN785
0T=?>YFgY]^[[OYa0=_MK5GKc528;,E+DHU@Cf1[B6I]R/:M&\QRW@1F/RR.ZSYY
8+RH>c,N=-S,YF0[O3X]CJ)=QB^D]O;DLM3:(P?5OdXM6WH[^W=Z+1_+b7UTBFPP
VJ3@YLVa>X/XGA_YbI[S(ODPNL(gRWMd1@^2T5\:8]/FC3<1:8QRZ1&ad<VZ31W9
6EK:>Kb1,-_gVC-^b>eJI:VASO_5ZJL/fTg[eY#X,BA?[;BV^TW,W\6XEddI1efK
fO5FZaNUPD1ANI.Z1eL6IVV/f;.[N@/ZT/5&1M.aXRa<./f6)]3I1^C\MYP)>\7e
M31NWTB:AF<,#72I,<LHDfY89?-6AaZZ;R@/^c)R#Sb:4b^\eR;,KegGH<(=>=YT
U_N0]c<H=J>LUa-0S#-9=[H2Bc0P-/Z[<\@NARa/>;QC6R=?XA&=G7BF.dX8J,E(
TWI2PMb+\+R3.S9+IKN0_L7J<?S?;CVRRRH38^[J:TH)[1\4Rbd@/MN450N)C-;(
DQ@PeBS<=If[\1@SF(0473=f3,6+AL^_]V<@be&;>_H)+f=BQX7fc#SFF1[;>^XN
PggcE/>Z79:8OTO[L9-)64gbB1()YY47:V0cE&.EcJ8_8UAGL>RZI?C#M?.KTd8=
=^-A?&c.2:[0U^=9HV_U2NfEKQS0)Bbf9R3;[8>OFR,+Q/bfX)HA9dCad47B-LW2
RGAcaLFV=8=LEf^cJ#VS8YU96/8<[-I5DKWU:D8-ZZ(]-QJ-]g=6bNaMS&9:16RS
G@-&]ea2[&B/RdD@J+K)W.0I[>I?P1c3g>3\L]J]FPK@+Q\Eebf5=Z0KX;U6F?:V
d\I6:c;3)6-;9;bPHZPMX:66KT+g^IVf9agDcI5IGS;PR,IMD)5)gVEced&W.cLa
QMHTSe8]BIO1Zf,76V-UOCS)33gR(XWe-1b^6HQQBg-DQ5JNKcPD=;DS(V:.3g&-
P4#/U1SFF(__W8BB]L-.ZP,.J-,?]MA<_cgAQ6fgLf70cS9^,38:ZMe\]<beN;5Q
H.@X;gQf1>8a[ULW(AFOaL3.&Oaa#\T?eJGd<]KBed@T:&baETb69f6>Kdg<)_R@
5fT@CT-OMg@c1QMKBg:S<W_0c;gK0^X>V:Q,4)Q989fBX4O6IY_)4YG+7/>(OD-Z
:5@NQIXBSOP4L=T&C+O(-TQ5ZfW9#/:g>&KN,JYS,[4gFacH4Q1L.dUbdYVSfIQA
f,J;,F\4<+a,NY]\IRYS]B^(Y5#8[RGgQgK/#?8X=>fQAfG0YfXJdddS=Q457R@,
P^,Qcf80gE>=216CAc:I&=:K7A&8Oc+KE/U0f9JIPPgIIMT-gHIR])bc.^T[gN\6
CcgU==57R;M#SE4\RE3G;D;bg)?<(BaP5+0Vba#LSb\3<#UDIX>:QRE3O+gMH7g&
:;41EX1DC?>#UNa8\6GeBYT3Z[O0U;I]2FT(@.1<A:P7;&PWEPYZV3H\]aIXNXbK
De7LY=:2C=5?]^I/SJ?9((RIAc\N[b_)/4FOB=D7QcJ3.&6QLEN>IF;YZ+[5@)L[
SUTVc8eV)RR=#]#7A,=JbL@.Y6M@3&8:_?=.C-gfYGeU@CgLZ1BZZO?bNUAb1NJ0
d;0XafXWU0;O;4:WW3B#9>N.^9?dL@[(1=HNKL7b-f&<TdQKVR&MZ9\0f&^cF\O-
Rb.<@FQ=S5;>S1c23.bR0K>7D[[fDU4[-\fF;)-KJ7\EFG5)(&g-<<f583UXT6E@
&S<97dI\W&S9>X1CU<(0&\?WNg.2b[LJQWUa<J1<BT0A6bPedeDFHH3T44E?75-]
_&>6W3<IOLQ9Sa14W5:V8TC29=@^KTd]YNfYBPN.JZc7OYbecG;K6@0IEdTTL@SF
P;23XSdB#[&]@YK3g+?/&00?QL__X>HRS5LSWRF4EM/B)2DbRGF]I1O^^]_A,]T@
dZ::?0g@&?V[Se?;_+WC=E?_X.<[LHgJ90TWC=:N#^K&H&]Y_QH_>RD6V,81HgF_
-dH^>,M_ScQ[C#2c&.830<3CgYA=9\K&=8ZKVWY7>5].&MOBQY4FYf66?CR8-cOF
=Ff>=dcU8LCFIb,(/3#J2[:3RL6K_:RgL-f;4P.dM#Y^g+3AJ>7E1I^^^Q^Q/64+
Q]RH&)#>&0^_C?]RD-B=[>Db@;LX,^egXZFB5H/KaA=31RQ.YgXQ857R8DZ4(DX@
RHF:)S,9>PS/CRIVe?O?A-3=R>OW[b;0fE=9\_S;DQL4d#[1FJ827=D#cPO\<RZ,
0D94=5cPOJ/=A2ZHN>PHP@@2A,1\Ef=IO[+a_/c5/e=]WZ@FP.B;GA-=ZFH5P+R/
-+JQ2F/aT:;86LIV2NB/(MO.FAON@#X_O>:XJ;^7/bT;TRD[1(>Rc2)D8FBcgb;X
ODSfBa3/ae=+?Ma/S[c0]b.V9DOE>6HAO925:8f&YJNV<5T0YB/O?11gd0gD(U:W
\_7[dc5V&_O:HE8,(1-d/5JNPW]-A(YSeCZJI8fe9&/7<b]),O5T>;91GbB5f5S1
FL[YYA+OENf=3O9TROB2-;/Y3DdSMZ\03&CEdIV.),.1Z;?Ff#4M2IfSH8c.F6NX
_Sed/7Z6H^.PPM79@@;YbYNQ8Q2Xc,YOS2f=@\Ngb86eJ^9NPT,SgV9Z;^U5EHTQ
O?X0T[AF1GHEGSGAK]59?#BT,];YY)S)V/e]JIfG9/7cN8dfVIH311AUQ1;Y_<<G
0f_OQHVQ83-)4.F3NP.UF6B4;aE7<4CJ,eYL\3(:YESK3C#1aNDV759EAbd8L;(P
K[6ff<DG8JYgf7UGBUMdOTP_b0gI63,?Tf00V[7+@UYF/g3DCPSBb1IM>S=eZ;6K
4#.J5(+8EZ-]N<\e@SQW@:>9Uf(UeeC7R8,];#-O0S#^?A#\JDO:N_8,,OOUX_ZQ
HIT],00/:K2^5WK/1=WZ:9.K59Y566?;f?73(KdZ5=R[bJbd^?X-C8\?XDA^MI\6
>:6F]Pefe715S96<cXBS(KRXM]>KJgLODBL?1JO\85=Tc.J4dD<:/Ebc^P1THc(C
[8X7F>LfV?dWOR7TVRP:9^T9]JF#a5]W[IB:V;-3SU6VJ6KOCb>S:BOR8M1L(8-L
G5VHH?.M;IP4[bBHR\?YKe0c3VSM;R@P^C;<-8_9L]I3TK4J=fSC@=5OQKZSD,N5
-gWORGg7P0K,]@;>YB1=N8dKJYZecGP;Uf/WO2aCPH[6ZQGO2BdCZZ.CP9d=&^>-
1Z&,Pb(P#IQfKN?Q2HW-^]1Pa-IE#X^J6SNII-V3<B,4O.S?#-+;1?3?4?M18WSc
L@6+EGKBLW3B:AZY?#W+R=.B\Id3g&RA?NZ&S)I^I<X72.[7;(,#SE#@A/e([]K<
d76YH==O[1cM.LLG2MGJOL>\]fDMB<KCQ#KJ\WU>b@NGV88V4JY5^?-dKV?#dGPQ
UG-Y090cF.(T<A(IDc<]@fW&)a#>7G5.7S1I^)/<aJ[L3;WBO,/28X4AZM\20b9J
O[0)5-JS>,-g=KTW)1f1)E7QUL7IK34J:#>YBNI).RF?<KC<e]g4_?FDXG1LQW<2
D\/Y]EA_81Ng&TK>8/+B+TH,(@>B4ZQE?LFZ@c=L8DZcT9LeTC@fFdCgRdMVKc=M
-CJ]e;:Q3V8K#,Y]FSZSAN-5cUX@aMa#+PK9NbG63W#/__+-8=fFad\(-\@F&.3:
K/fBSM4PcYMKXM4[d\^^caB&[(IdO<Nb+b_YXK-Y+6HZN9UEbXNTALEf3].];.3L
<4e)774/Qb\;<G1QQcAc^-J4Y(?43[K7f(A-aAd#.RSY1Ve+HBS@K(1I78D>>V&A
1e?5>U0Bf#IJ05?C;@6N_6]NT)C9>a-_Q\gS;BF0d.)fP[--)O>8NP43<HR:ee^d
P\AL281eN_KZ671a,P4dcTG_PM]cb2>YcIU^)9f0F_^eEATQCHcfe+W)DHIN5OUO
V1&A/KOTLLO;,<HgdALgPdYVVCHPR/EA6WM[[-J#Z6HDR5L1\RP/W>GB(EA>ZR]^
Oc\/<XKVN[eLA#?O/aO25H1(aSJ_&5Q_c8BXPCHQT36UT7[=0=a6dc[bWJ^cGJ_M
HSebbNPdQ#R&BA+aV9T>[5aM/Y8+U</0J_bD?LWJLcA,aKCL&a\+6g,PKFEBb/,Y
U>E8f8Z@VE#:SQTBc-E5Q<J-8OBCBfg6D^gLb<>(dGNeT>]&VKB9O4+aFJU2[\JO
VB9c.NF?b/K2eD(=;aU[g4S>cJ<OI/\+94Y&,cRbJPA?caIH@5^])]N651Re5#[C
:P3ANP5/fJ8E^]QP1;ZV<;d/A25fgU853FKU(bZgRP>(,VJ&?2LR,K87e?RaK;?Z
#+1:6EAaH08M6HK^8TV725R9YHaW;fQH6E?^6(_BIC\PBTW399WCDHPfSEU\YG^a
5fJaJ5O&H-\>-[#EGWbOe<c0VY1?E7PeXSf/S[SO]@DM&.:@)ZG,::3\e<;3=RaX
.1dJRIG(g?[WbK.d5:)1,.HWa9BQ6)?J65-DH2D>Ma=@d7g59&,QUT]B8U03)FO5
L.f&K[^E:JdF93SRR&PV4#TaM:[>@)<JD=?;G^+-+C^_3M\(:YZQYWe3-EVGIWBR
d]Z:SOa5@ANJ0EV1Wa5-?OaY)@R3F2\Q,].=#_(F1baX,#;]ceZa?4AK(B\83b\K
BJ-g<S<=:f:?Gg3L1cUa5+<I@N)62I7e4f?@XbFHDGc6F\<Y-99M,g/fHQ064f3&
\6ZQD;J2K6BQ]<@/cF)OD#cf&&DM;/P>FAZCX,KP4U/MF+ed9)bOD@U?\E57JQ66
/:)f\@64EYK\HB1KD&bC&(WcFP3b_55f(R3ZH1#9B@aO3FgdeOOdV]eQ_a1350Xf
LB+I:C<V[1REE[?+0G1OQg:]FHY=;Z1)4fC&CX8[]Pd]G>L+.&V-/\PF\Bc4=NNe
1X<)];53I@()5(&P:((a-(1d3_M&RN>VG,P;9?&-@BY_LK+>cEH5K&4DYZD#9ZQD
?QF,,N=Fc3+78<f.UB>8fbNUHJJL+<Oa.#9K?_d;V;;HgSVJ]&fNIDf/FZ^a15>G
972AE6SU:UQ+G5=dKT9_dVdW?4C,Q&,8T\)P<+ZR\3?Pd+[:1AXWgHB65^eY)7N/
,dT#Z,9FH7>^RXRf@KV&eC6?\f=#BbV9(SR42f[bT]GRZMCX=GeFe+cV]:TD_5H6
K]gUC.A/)D\AX@Q:G)C-79;^\1##4aAZCMPB&?L7CZV;aR<BYS,NC-T4QWKd-V@>
04I-VNMcWV[[g^Z^-HVGCAA5<)Vbg8L[0e_.]65;9-K(#3PeE-4FP,Z[DSRKJCcA
RZ_TNQQ-@7P2^N_gV=e?<TgQ&__4AI-@M3(T8&K<#2gAfcH,D2Z83WBeQ@&I@2H^
VP]+cHO]]C&?OJd,0-E?]),#H4Y4+f.e2e#GKF--H+@S)/JUORbcB)BAI1_6F<BF
^FY3.=CS\O5)=]c]XfGTg7IeHM;-)RF5P7.1W)5/YCZ_E2AR8S39Mc).eK/>Q44f
-[GG<b]&V,(>1D7<fc&>-.RS+(;K<b2L+SS:(G;A&bBVaH@-8fK]_QGO:WgPJYP=
_+L].YcABfB)E1a;B[dPLaS,LFQEJ[>_?Y0[XTYCc;fDER2a>(X#:+=D9YLVdURH
SOb2ZdJ+WccC;b<=DHa+R1)]Ab9QXLTeMBP6e=^d&P<.YbdN?QQ&;?)UA:36:7gJ
_J;QHUa?)OYYWCQBQDU=?#AZZc0C<P-T/U9XB=-LVO?CMIZfQF3SJNSIF-dYZ@=Q
b;YCeNO?D-BSc;faT5NG6CcV:26<[aHFE=fY7bfOWeLVW-3GUF>@.,YfQND-63#I
TB58.?COFV=V8-===<KCN)4IGL<<?@I3=EQ39_b^:1R)e2C,dVRT2H/UGf0]cdD5
Q=I:B/a;V7NZI[0#^^:2e0VdM<KN:.L1,S^,A))SOIM,\)-QA\><D;f1;EP:#O[f
adX_;JIZ+Ja=9_C).SKPXb7>=L,2Q+8BA]V-T<<BGC[48d-]-RN^^?bT5?C#6(cR
.d;C<T+M.T1,YbaM&DE.<(,+F.U[SVe@02fPAAB\B(X:a>^Z&T]4TQ<8X)^6=,?]
Q5\4,?Q1f:_gKDb^17g;[GNLFM&fL8M^WG[<I0ND8cDc?Ue,F0@SQ?RS[,O1,/7E
T9T5S=VJU#+&H^2c14NT154R[(X&2+QLceCHB4FaC>b65.caU\BSOdPHA#Kdge.4
PSMAXP9:VB,ON\CWZ;LY_1QJ5-c9S-)DNLH?,Z^1;7[^#>9/1RSeC-aRZNPQU:N1
51R4c.SLcPP(Hg2[&C;QK@D;^b<BGbb/)Bg=H.;).>Z?D]UE+6_e<&K^B&\KRGdK
7N3/9LZZ;=PN:4^<RT[8/Ug[E0E>d\W+/)\_:dg.E&dE9EZS?_):bI0EFg7&#[KA
cTH4GD;@g.TM1X^Z-I9^_a,aAeA-7@:5U=XSLPENdHg[(I4BPg>d##A:F94]_Y?;
5:36U4])O??.#HeGXWc1=AJR4[ZS9cc,:@((4,[>G+H/K-ceWFN:E-HS=5-B<I<E
IHL];,NdARFL=;R)f<]Z@]2TJ/13[B742Z3f75[BeN@3BZ6:^2O5;4V_c3+EEN-P
^c)7[cL33@XP?U9F8E:f[^f4)VIb]\)2]ZOP]@<\]G)5g[UO5cI70]YIKd.T6L[J
0IC5XaYXgUW?1eLfX)+IC7+1,S2#1MFJ0Ag/#\Re>MMA-Q-#d&^+NQ,3agK(,>3f
AYE7.68;;CC,_VLAZS6+gET\PWA2>&,ACQaG-R^M6K>P)AXD>0?(<g(T[7Na?4>J
::6AV]SZ,P8&5;8/&A0]6dK&>Z+PL_fJIMZ/&<L[@=U+XfG=.Q9/XA&UXZ=E[U2<
VV]WJC4.CM^.#&#:Na=UPVd=KAH4G5DA8efXNVQW6EC-bf^]A7fRJV0/7D<KUf_1
;1H2UaSJSO0[,M,X.#(HX+-HI]P)/Y^BLR2=GI&P?,bULa>-,.38C5OK4XMW=G:4
d?:IEL^?d9N;NVGg#9JC2A)BJMGQBF1<Z7J-gd0X<(Ab[5ZNf2#K_\6Q_^>7#J\L
.X56,,-eK]./TFS1NcDT/-Z8>@M)LF#HSGB2].<)8_X:Z(W[?]f6?\DS/G()5,gB
a>D)E01U.+F/17a8JF)KIKK<[1b?@)F,+QB14EeO_TFUd3G]]:_W)=@&66c)].O5
7e5Q(_&.J1++/4_\1)AH.EP;b@[Y4T-;UZ&=d;#>Z?1&XMT+bgUaSC_PD090.6ea
9;W8BD(1ZJ>B]:)9VV4=9RA:+9M>B0^P^1JH.X2/DZ&(EF10I#;ag=+LI;0d[2Oc
VNI^,O7BA-/b<]27EDH,4JK-Sa/7Vc,Y3-Te8^>79/fFX&HNOG3Bd(;c0T>W+8ZC
f60fdNHP2J/:cQ)HBM3gJGHJG0AU997PKE8a-=#@2H.A]X:6aI8(SC@Me)FbI\BR
T[\YgBRB=AB[bId7.;GWIK&,].4F:::bdZ<35C(LRXc>dCV<B&P)(QI/;IHO>dcN
52UNJ=DD\D,:gDZ[CQ??LGgb(f]Bf^/a5JXcR1NPZ3QYZF_2X@R_6f\JRGO7H8Q4
K34]N5YC>.T.Pa=GS8&c3@\(V#S[E;EDg(77D4J_BJK_M9\;>/#M)SDg=/+5&a/V
U@FHEG(3bR8SX7_C.6dF@4QI<)+7A<8I16B1g#8(IM-&RUc+S=_F@8(ZR?OBK2\Y
5IXZgB(5DTX-OCQff@1-D]T8BfYZJ)._W@a?A1-_?,]TUS_D1_8?87K<?NY.\&AX
:eP==24_-a+MJ(fcY)2CYEKO79F,6&]JKGNV9SRAGMNa\6f.HPa76C@Xc&:MY)fI
c/[5^#PdeYB6;5AFE7F,9SKO2$
`endprotected
endmodule


