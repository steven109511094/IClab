# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : mem_ker
#       Words            : 80
#       Bits             : 40
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/03/29 20:04:00
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO mem_ker
CLASS BLOCK ;
FOREIGN mem_ker 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 655.340 BY 161.840 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 654.220 129.700 655.340 132.940 ;
  LAYER ME3 ;
  RECT 654.220 129.700 655.340 132.940 ;
  LAYER ME2 ;
  RECT 654.220 129.700 655.340 132.940 ;
  LAYER ME1 ;
  RECT 654.220 129.700 655.340 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 121.860 655.340 125.100 ;
  LAYER ME3 ;
  RECT 654.220 121.860 655.340 125.100 ;
  LAYER ME2 ;
  RECT 654.220 121.860 655.340 125.100 ;
  LAYER ME1 ;
  RECT 654.220 121.860 655.340 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 114.020 655.340 117.260 ;
  LAYER ME3 ;
  RECT 654.220 114.020 655.340 117.260 ;
  LAYER ME2 ;
  RECT 654.220 114.020 655.340 117.260 ;
  LAYER ME1 ;
  RECT 654.220 114.020 655.340 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 106.180 655.340 109.420 ;
  LAYER ME3 ;
  RECT 654.220 106.180 655.340 109.420 ;
  LAYER ME2 ;
  RECT 654.220 106.180 655.340 109.420 ;
  LAYER ME1 ;
  RECT 654.220 106.180 655.340 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 98.340 655.340 101.580 ;
  LAYER ME3 ;
  RECT 654.220 98.340 655.340 101.580 ;
  LAYER ME2 ;
  RECT 654.220 98.340 655.340 101.580 ;
  LAYER ME1 ;
  RECT 654.220 98.340 655.340 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 90.500 655.340 93.740 ;
  LAYER ME3 ;
  RECT 654.220 90.500 655.340 93.740 ;
  LAYER ME2 ;
  RECT 654.220 90.500 655.340 93.740 ;
  LAYER ME1 ;
  RECT 654.220 90.500 655.340 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 51.300 655.340 54.540 ;
  LAYER ME3 ;
  RECT 654.220 51.300 655.340 54.540 ;
  LAYER ME2 ;
  RECT 654.220 51.300 655.340 54.540 ;
  LAYER ME1 ;
  RECT 654.220 51.300 655.340 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 43.460 655.340 46.700 ;
  LAYER ME3 ;
  RECT 654.220 43.460 655.340 46.700 ;
  LAYER ME2 ;
  RECT 654.220 43.460 655.340 46.700 ;
  LAYER ME1 ;
  RECT 654.220 43.460 655.340 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 35.620 655.340 38.860 ;
  LAYER ME3 ;
  RECT 654.220 35.620 655.340 38.860 ;
  LAYER ME2 ;
  RECT 654.220 35.620 655.340 38.860 ;
  LAYER ME1 ;
  RECT 654.220 35.620 655.340 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 27.780 655.340 31.020 ;
  LAYER ME3 ;
  RECT 654.220 27.780 655.340 31.020 ;
  LAYER ME2 ;
  RECT 654.220 27.780 655.340 31.020 ;
  LAYER ME1 ;
  RECT 654.220 27.780 655.340 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 19.940 655.340 23.180 ;
  LAYER ME3 ;
  RECT 654.220 19.940 655.340 23.180 ;
  LAYER ME2 ;
  RECT 654.220 19.940 655.340 23.180 ;
  LAYER ME1 ;
  RECT 654.220 19.940 655.340 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 12.100 655.340 15.340 ;
  LAYER ME3 ;
  RECT 654.220 12.100 655.340 15.340 ;
  LAYER ME2 ;
  RECT 654.220 12.100 655.340 15.340 ;
  LAYER ME1 ;
  RECT 654.220 12.100 655.340 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 637.140 160.720 640.680 161.840 ;
  LAYER ME3 ;
  RECT 637.140 160.720 640.680 161.840 ;
  LAYER ME2 ;
  RECT 637.140 160.720 640.680 161.840 ;
  LAYER ME1 ;
  RECT 637.140 160.720 640.680 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 628.460 160.720 632.000 161.840 ;
  LAYER ME3 ;
  RECT 628.460 160.720 632.000 161.840 ;
  LAYER ME2 ;
  RECT 628.460 160.720 632.000 161.840 ;
  LAYER ME1 ;
  RECT 628.460 160.720 632.000 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 619.780 160.720 623.320 161.840 ;
  LAYER ME3 ;
  RECT 619.780 160.720 623.320 161.840 ;
  LAYER ME2 ;
  RECT 619.780 160.720 623.320 161.840 ;
  LAYER ME1 ;
  RECT 619.780 160.720 623.320 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 576.380 160.720 579.920 161.840 ;
  LAYER ME3 ;
  RECT 576.380 160.720 579.920 161.840 ;
  LAYER ME2 ;
  RECT 576.380 160.720 579.920 161.840 ;
  LAYER ME1 ;
  RECT 576.380 160.720 579.920 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 567.700 160.720 571.240 161.840 ;
  LAYER ME3 ;
  RECT 567.700 160.720 571.240 161.840 ;
  LAYER ME2 ;
  RECT 567.700 160.720 571.240 161.840 ;
  LAYER ME1 ;
  RECT 567.700 160.720 571.240 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 559.020 160.720 562.560 161.840 ;
  LAYER ME3 ;
  RECT 559.020 160.720 562.560 161.840 ;
  LAYER ME2 ;
  RECT 559.020 160.720 562.560 161.840 ;
  LAYER ME1 ;
  RECT 559.020 160.720 562.560 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 550.340 160.720 553.880 161.840 ;
  LAYER ME3 ;
  RECT 550.340 160.720 553.880 161.840 ;
  LAYER ME2 ;
  RECT 550.340 160.720 553.880 161.840 ;
  LAYER ME1 ;
  RECT 550.340 160.720 553.880 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 541.660 160.720 545.200 161.840 ;
  LAYER ME3 ;
  RECT 541.660 160.720 545.200 161.840 ;
  LAYER ME2 ;
  RECT 541.660 160.720 545.200 161.840 ;
  LAYER ME1 ;
  RECT 541.660 160.720 545.200 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 532.980 160.720 536.520 161.840 ;
  LAYER ME3 ;
  RECT 532.980 160.720 536.520 161.840 ;
  LAYER ME2 ;
  RECT 532.980 160.720 536.520 161.840 ;
  LAYER ME1 ;
  RECT 532.980 160.720 536.520 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 160.720 493.120 161.840 ;
  LAYER ME3 ;
  RECT 489.580 160.720 493.120 161.840 ;
  LAYER ME2 ;
  RECT 489.580 160.720 493.120 161.840 ;
  LAYER ME1 ;
  RECT 489.580 160.720 493.120 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 160.720 484.440 161.840 ;
  LAYER ME3 ;
  RECT 480.900 160.720 484.440 161.840 ;
  LAYER ME2 ;
  RECT 480.900 160.720 484.440 161.840 ;
  LAYER ME1 ;
  RECT 480.900 160.720 484.440 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 160.720 475.760 161.840 ;
  LAYER ME3 ;
  RECT 472.220 160.720 475.760 161.840 ;
  LAYER ME2 ;
  RECT 472.220 160.720 475.760 161.840 ;
  LAYER ME1 ;
  RECT 472.220 160.720 475.760 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 160.720 467.080 161.840 ;
  LAYER ME3 ;
  RECT 463.540 160.720 467.080 161.840 ;
  LAYER ME2 ;
  RECT 463.540 160.720 467.080 161.840 ;
  LAYER ME1 ;
  RECT 463.540 160.720 467.080 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 160.720 458.400 161.840 ;
  LAYER ME3 ;
  RECT 454.860 160.720 458.400 161.840 ;
  LAYER ME2 ;
  RECT 454.860 160.720 458.400 161.840 ;
  LAYER ME1 ;
  RECT 454.860 160.720 458.400 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 160.720 449.720 161.840 ;
  LAYER ME3 ;
  RECT 446.180 160.720 449.720 161.840 ;
  LAYER ME2 ;
  RECT 446.180 160.720 449.720 161.840 ;
  LAYER ME1 ;
  RECT 446.180 160.720 449.720 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 160.720 406.320 161.840 ;
  LAYER ME3 ;
  RECT 402.780 160.720 406.320 161.840 ;
  LAYER ME2 ;
  RECT 402.780 160.720 406.320 161.840 ;
  LAYER ME1 ;
  RECT 402.780 160.720 406.320 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 160.720 397.640 161.840 ;
  LAYER ME3 ;
  RECT 394.100 160.720 397.640 161.840 ;
  LAYER ME2 ;
  RECT 394.100 160.720 397.640 161.840 ;
  LAYER ME1 ;
  RECT 394.100 160.720 397.640 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 160.720 388.960 161.840 ;
  LAYER ME3 ;
  RECT 385.420 160.720 388.960 161.840 ;
  LAYER ME2 ;
  RECT 385.420 160.720 388.960 161.840 ;
  LAYER ME1 ;
  RECT 385.420 160.720 388.960 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 160.720 380.280 161.840 ;
  LAYER ME3 ;
  RECT 376.740 160.720 380.280 161.840 ;
  LAYER ME2 ;
  RECT 376.740 160.720 380.280 161.840 ;
  LAYER ME1 ;
  RECT 376.740 160.720 380.280 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 160.720 371.600 161.840 ;
  LAYER ME3 ;
  RECT 368.060 160.720 371.600 161.840 ;
  LAYER ME2 ;
  RECT 368.060 160.720 371.600 161.840 ;
  LAYER ME1 ;
  RECT 368.060 160.720 371.600 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 160.720 362.920 161.840 ;
  LAYER ME3 ;
  RECT 359.380 160.720 362.920 161.840 ;
  LAYER ME2 ;
  RECT 359.380 160.720 362.920 161.840 ;
  LAYER ME1 ;
  RECT 359.380 160.720 362.920 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 160.720 319.520 161.840 ;
  LAYER ME3 ;
  RECT 315.980 160.720 319.520 161.840 ;
  LAYER ME2 ;
  RECT 315.980 160.720 319.520 161.840 ;
  LAYER ME1 ;
  RECT 315.980 160.720 319.520 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 160.720 310.840 161.840 ;
  LAYER ME3 ;
  RECT 307.300 160.720 310.840 161.840 ;
  LAYER ME2 ;
  RECT 307.300 160.720 310.840 161.840 ;
  LAYER ME1 ;
  RECT 307.300 160.720 310.840 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 160.720 302.160 161.840 ;
  LAYER ME3 ;
  RECT 298.620 160.720 302.160 161.840 ;
  LAYER ME2 ;
  RECT 298.620 160.720 302.160 161.840 ;
  LAYER ME1 ;
  RECT 298.620 160.720 302.160 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 160.720 293.480 161.840 ;
  LAYER ME3 ;
  RECT 289.940 160.720 293.480 161.840 ;
  LAYER ME2 ;
  RECT 289.940 160.720 293.480 161.840 ;
  LAYER ME1 ;
  RECT 289.940 160.720 293.480 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 160.720 284.800 161.840 ;
  LAYER ME3 ;
  RECT 281.260 160.720 284.800 161.840 ;
  LAYER ME2 ;
  RECT 281.260 160.720 284.800 161.840 ;
  LAYER ME1 ;
  RECT 281.260 160.720 284.800 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 160.720 276.120 161.840 ;
  LAYER ME3 ;
  RECT 272.580 160.720 276.120 161.840 ;
  LAYER ME2 ;
  RECT 272.580 160.720 276.120 161.840 ;
  LAYER ME1 ;
  RECT 272.580 160.720 276.120 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 160.720 232.720 161.840 ;
  LAYER ME3 ;
  RECT 229.180 160.720 232.720 161.840 ;
  LAYER ME2 ;
  RECT 229.180 160.720 232.720 161.840 ;
  LAYER ME1 ;
  RECT 229.180 160.720 232.720 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 160.720 224.040 161.840 ;
  LAYER ME3 ;
  RECT 220.500 160.720 224.040 161.840 ;
  LAYER ME2 ;
  RECT 220.500 160.720 224.040 161.840 ;
  LAYER ME1 ;
  RECT 220.500 160.720 224.040 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 160.720 215.360 161.840 ;
  LAYER ME3 ;
  RECT 211.820 160.720 215.360 161.840 ;
  LAYER ME2 ;
  RECT 211.820 160.720 215.360 161.840 ;
  LAYER ME1 ;
  RECT 211.820 160.720 215.360 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 160.720 206.680 161.840 ;
  LAYER ME3 ;
  RECT 203.140 160.720 206.680 161.840 ;
  LAYER ME2 ;
  RECT 203.140 160.720 206.680 161.840 ;
  LAYER ME1 ;
  RECT 203.140 160.720 206.680 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 160.720 198.000 161.840 ;
  LAYER ME3 ;
  RECT 194.460 160.720 198.000 161.840 ;
  LAYER ME2 ;
  RECT 194.460 160.720 198.000 161.840 ;
  LAYER ME1 ;
  RECT 194.460 160.720 198.000 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 160.720 189.320 161.840 ;
  LAYER ME3 ;
  RECT 185.780 160.720 189.320 161.840 ;
  LAYER ME2 ;
  RECT 185.780 160.720 189.320 161.840 ;
  LAYER ME1 ;
  RECT 185.780 160.720 189.320 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 160.720 145.920 161.840 ;
  LAYER ME3 ;
  RECT 142.380 160.720 145.920 161.840 ;
  LAYER ME2 ;
  RECT 142.380 160.720 145.920 161.840 ;
  LAYER ME1 ;
  RECT 142.380 160.720 145.920 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 160.720 137.240 161.840 ;
  LAYER ME3 ;
  RECT 133.700 160.720 137.240 161.840 ;
  LAYER ME2 ;
  RECT 133.700 160.720 137.240 161.840 ;
  LAYER ME1 ;
  RECT 133.700 160.720 137.240 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 160.720 128.560 161.840 ;
  LAYER ME3 ;
  RECT 125.020 160.720 128.560 161.840 ;
  LAYER ME2 ;
  RECT 125.020 160.720 128.560 161.840 ;
  LAYER ME1 ;
  RECT 125.020 160.720 128.560 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 160.720 119.880 161.840 ;
  LAYER ME3 ;
  RECT 116.340 160.720 119.880 161.840 ;
  LAYER ME2 ;
  RECT 116.340 160.720 119.880 161.840 ;
  LAYER ME1 ;
  RECT 116.340 160.720 119.880 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 160.720 111.200 161.840 ;
  LAYER ME3 ;
  RECT 107.660 160.720 111.200 161.840 ;
  LAYER ME2 ;
  RECT 107.660 160.720 111.200 161.840 ;
  LAYER ME1 ;
  RECT 107.660 160.720 111.200 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 160.720 102.520 161.840 ;
  LAYER ME3 ;
  RECT 98.980 160.720 102.520 161.840 ;
  LAYER ME2 ;
  RECT 98.980 160.720 102.520 161.840 ;
  LAYER ME1 ;
  RECT 98.980 160.720 102.520 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 160.720 59.120 161.840 ;
  LAYER ME3 ;
  RECT 55.580 160.720 59.120 161.840 ;
  LAYER ME2 ;
  RECT 55.580 160.720 59.120 161.840 ;
  LAYER ME1 ;
  RECT 55.580 160.720 59.120 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 160.720 50.440 161.840 ;
  LAYER ME3 ;
  RECT 46.900 160.720 50.440 161.840 ;
  LAYER ME2 ;
  RECT 46.900 160.720 50.440 161.840 ;
  LAYER ME1 ;
  RECT 46.900 160.720 50.440 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 160.720 41.760 161.840 ;
  LAYER ME3 ;
  RECT 38.220 160.720 41.760 161.840 ;
  LAYER ME2 ;
  RECT 38.220 160.720 41.760 161.840 ;
  LAYER ME1 ;
  RECT 38.220 160.720 41.760 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 160.720 33.080 161.840 ;
  LAYER ME3 ;
  RECT 29.540 160.720 33.080 161.840 ;
  LAYER ME2 ;
  RECT 29.540 160.720 33.080 161.840 ;
  LAYER ME1 ;
  RECT 29.540 160.720 33.080 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 160.720 24.400 161.840 ;
  LAYER ME3 ;
  RECT 20.860 160.720 24.400 161.840 ;
  LAYER ME2 ;
  RECT 20.860 160.720 24.400 161.840 ;
  LAYER ME1 ;
  RECT 20.860 160.720 24.400 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 160.720 15.720 161.840 ;
  LAYER ME3 ;
  RECT 12.180 160.720 15.720 161.840 ;
  LAYER ME2 ;
  RECT 12.180 160.720 15.720 161.840 ;
  LAYER ME1 ;
  RECT 12.180 160.720 15.720 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME3 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME2 ;
  RECT 565.840 0.000 569.380 1.120 ;
  LAYER ME1 ;
  RECT 565.840 0.000 569.380 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME3 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME2 ;
  RECT 549.100 0.000 552.640 1.120 ;
  LAYER ME1 ;
  RECT 549.100 0.000 552.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME3 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME2 ;
  RECT 522.440 0.000 525.980 1.120 ;
  LAYER ME1 ;
  RECT 522.440 0.000 525.980 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME3 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME2 ;
  RECT 500.740 0.000 504.280 1.120 ;
  LAYER ME1 ;
  RECT 500.740 0.000 504.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME3 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME2 ;
  RECT 479.660 0.000 483.200 1.120 ;
  LAYER ME1 ;
  RECT 479.660 0.000 483.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME3 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME2 ;
  RECT 453.000 0.000 456.540 1.120 ;
  LAYER ME1 ;
  RECT 453.000 0.000 456.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME3 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME2 ;
  RECT 339.540 0.000 343.080 1.120 ;
  LAYER ME1 ;
  RECT 339.540 0.000 343.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER ME3 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER ME2 ;
  RECT 330.860 0.000 334.400 1.120 ;
  LAYER ME1 ;
  RECT 330.860 0.000 334.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 0.000 306.500 1.120 ;
  LAYER ME3 ;
  RECT 302.960 0.000 306.500 1.120 ;
  LAYER ME2 ;
  RECT 302.960 0.000 306.500 1.120 ;
  LAYER ME1 ;
  RECT 302.960 0.000 306.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 291.800 0.000 295.340 1.120 ;
  LAYER ME3 ;
  RECT 291.800 0.000 295.340 1.120 ;
  LAYER ME2 ;
  RECT 291.800 0.000 295.340 1.120 ;
  LAYER ME1 ;
  RECT 291.800 0.000 295.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME3 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME2 ;
  RECT 270.100 0.000 273.640 1.120 ;
  LAYER ME1 ;
  RECT 270.100 0.000 273.640 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME3 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME2 ;
  RECT 253.360 0.000 256.900 1.120 ;
  LAYER ME1 ;
  RECT 253.360 0.000 256.900 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 654.220 125.780 655.340 129.020 ;
  LAYER ME3 ;
  RECT 654.220 125.780 655.340 129.020 ;
  LAYER ME2 ;
  RECT 654.220 125.780 655.340 129.020 ;
  LAYER ME1 ;
  RECT 654.220 125.780 655.340 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 117.940 655.340 121.180 ;
  LAYER ME3 ;
  RECT 654.220 117.940 655.340 121.180 ;
  LAYER ME2 ;
  RECT 654.220 117.940 655.340 121.180 ;
  LAYER ME1 ;
  RECT 654.220 117.940 655.340 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 110.100 655.340 113.340 ;
  LAYER ME3 ;
  RECT 654.220 110.100 655.340 113.340 ;
  LAYER ME2 ;
  RECT 654.220 110.100 655.340 113.340 ;
  LAYER ME1 ;
  RECT 654.220 110.100 655.340 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 102.260 655.340 105.500 ;
  LAYER ME3 ;
  RECT 654.220 102.260 655.340 105.500 ;
  LAYER ME2 ;
  RECT 654.220 102.260 655.340 105.500 ;
  LAYER ME1 ;
  RECT 654.220 102.260 655.340 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 94.420 655.340 97.660 ;
  LAYER ME3 ;
  RECT 654.220 94.420 655.340 97.660 ;
  LAYER ME2 ;
  RECT 654.220 94.420 655.340 97.660 ;
  LAYER ME1 ;
  RECT 654.220 94.420 655.340 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 86.580 655.340 89.820 ;
  LAYER ME3 ;
  RECT 654.220 86.580 655.340 89.820 ;
  LAYER ME2 ;
  RECT 654.220 86.580 655.340 89.820 ;
  LAYER ME1 ;
  RECT 654.220 86.580 655.340 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 47.380 655.340 50.620 ;
  LAYER ME3 ;
  RECT 654.220 47.380 655.340 50.620 ;
  LAYER ME2 ;
  RECT 654.220 47.380 655.340 50.620 ;
  LAYER ME1 ;
  RECT 654.220 47.380 655.340 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 39.540 655.340 42.780 ;
  LAYER ME3 ;
  RECT 654.220 39.540 655.340 42.780 ;
  LAYER ME2 ;
  RECT 654.220 39.540 655.340 42.780 ;
  LAYER ME1 ;
  RECT 654.220 39.540 655.340 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 31.700 655.340 34.940 ;
  LAYER ME3 ;
  RECT 654.220 31.700 655.340 34.940 ;
  LAYER ME2 ;
  RECT 654.220 31.700 655.340 34.940 ;
  LAYER ME1 ;
  RECT 654.220 31.700 655.340 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 23.860 655.340 27.100 ;
  LAYER ME3 ;
  RECT 654.220 23.860 655.340 27.100 ;
  LAYER ME2 ;
  RECT 654.220 23.860 655.340 27.100 ;
  LAYER ME1 ;
  RECT 654.220 23.860 655.340 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 16.020 655.340 19.260 ;
  LAYER ME3 ;
  RECT 654.220 16.020 655.340 19.260 ;
  LAYER ME2 ;
  RECT 654.220 16.020 655.340 19.260 ;
  LAYER ME1 ;
  RECT 654.220 16.020 655.340 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 654.220 8.180 655.340 11.420 ;
  LAYER ME3 ;
  RECT 654.220 8.180 655.340 11.420 ;
  LAYER ME2 ;
  RECT 654.220 8.180 655.340 11.420 ;
  LAYER ME1 ;
  RECT 654.220 8.180 655.340 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 641.480 160.720 645.020 161.840 ;
  LAYER ME3 ;
  RECT 641.480 160.720 645.020 161.840 ;
  LAYER ME2 ;
  RECT 641.480 160.720 645.020 161.840 ;
  LAYER ME1 ;
  RECT 641.480 160.720 645.020 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 632.800 160.720 636.340 161.840 ;
  LAYER ME3 ;
  RECT 632.800 160.720 636.340 161.840 ;
  LAYER ME2 ;
  RECT 632.800 160.720 636.340 161.840 ;
  LAYER ME1 ;
  RECT 632.800 160.720 636.340 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 624.120 160.720 627.660 161.840 ;
  LAYER ME3 ;
  RECT 624.120 160.720 627.660 161.840 ;
  LAYER ME2 ;
  RECT 624.120 160.720 627.660 161.840 ;
  LAYER ME1 ;
  RECT 624.120 160.720 627.660 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 615.440 160.720 618.980 161.840 ;
  LAYER ME3 ;
  RECT 615.440 160.720 618.980 161.840 ;
  LAYER ME2 ;
  RECT 615.440 160.720 618.980 161.840 ;
  LAYER ME1 ;
  RECT 615.440 160.720 618.980 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 572.040 160.720 575.580 161.840 ;
  LAYER ME3 ;
  RECT 572.040 160.720 575.580 161.840 ;
  LAYER ME2 ;
  RECT 572.040 160.720 575.580 161.840 ;
  LAYER ME1 ;
  RECT 572.040 160.720 575.580 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 563.360 160.720 566.900 161.840 ;
  LAYER ME3 ;
  RECT 563.360 160.720 566.900 161.840 ;
  LAYER ME2 ;
  RECT 563.360 160.720 566.900 161.840 ;
  LAYER ME1 ;
  RECT 563.360 160.720 566.900 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 554.680 160.720 558.220 161.840 ;
  LAYER ME3 ;
  RECT 554.680 160.720 558.220 161.840 ;
  LAYER ME2 ;
  RECT 554.680 160.720 558.220 161.840 ;
  LAYER ME1 ;
  RECT 554.680 160.720 558.220 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 546.000 160.720 549.540 161.840 ;
  LAYER ME3 ;
  RECT 546.000 160.720 549.540 161.840 ;
  LAYER ME2 ;
  RECT 546.000 160.720 549.540 161.840 ;
  LAYER ME1 ;
  RECT 546.000 160.720 549.540 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 537.320 160.720 540.860 161.840 ;
  LAYER ME3 ;
  RECT 537.320 160.720 540.860 161.840 ;
  LAYER ME2 ;
  RECT 537.320 160.720 540.860 161.840 ;
  LAYER ME1 ;
  RECT 537.320 160.720 540.860 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 528.640 160.720 532.180 161.840 ;
  LAYER ME3 ;
  RECT 528.640 160.720 532.180 161.840 ;
  LAYER ME2 ;
  RECT 528.640 160.720 532.180 161.840 ;
  LAYER ME1 ;
  RECT 528.640 160.720 532.180 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 160.720 488.780 161.840 ;
  LAYER ME3 ;
  RECT 485.240 160.720 488.780 161.840 ;
  LAYER ME2 ;
  RECT 485.240 160.720 488.780 161.840 ;
  LAYER ME1 ;
  RECT 485.240 160.720 488.780 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 160.720 480.100 161.840 ;
  LAYER ME3 ;
  RECT 476.560 160.720 480.100 161.840 ;
  LAYER ME2 ;
  RECT 476.560 160.720 480.100 161.840 ;
  LAYER ME1 ;
  RECT 476.560 160.720 480.100 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 160.720 471.420 161.840 ;
  LAYER ME3 ;
  RECT 467.880 160.720 471.420 161.840 ;
  LAYER ME2 ;
  RECT 467.880 160.720 471.420 161.840 ;
  LAYER ME1 ;
  RECT 467.880 160.720 471.420 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 160.720 462.740 161.840 ;
  LAYER ME3 ;
  RECT 459.200 160.720 462.740 161.840 ;
  LAYER ME2 ;
  RECT 459.200 160.720 462.740 161.840 ;
  LAYER ME1 ;
  RECT 459.200 160.720 462.740 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 160.720 454.060 161.840 ;
  LAYER ME3 ;
  RECT 450.520 160.720 454.060 161.840 ;
  LAYER ME2 ;
  RECT 450.520 160.720 454.060 161.840 ;
  LAYER ME1 ;
  RECT 450.520 160.720 454.060 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 160.720 445.380 161.840 ;
  LAYER ME3 ;
  RECT 441.840 160.720 445.380 161.840 ;
  LAYER ME2 ;
  RECT 441.840 160.720 445.380 161.840 ;
  LAYER ME1 ;
  RECT 441.840 160.720 445.380 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 160.720 401.980 161.840 ;
  LAYER ME3 ;
  RECT 398.440 160.720 401.980 161.840 ;
  LAYER ME2 ;
  RECT 398.440 160.720 401.980 161.840 ;
  LAYER ME1 ;
  RECT 398.440 160.720 401.980 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 160.720 393.300 161.840 ;
  LAYER ME3 ;
  RECT 389.760 160.720 393.300 161.840 ;
  LAYER ME2 ;
  RECT 389.760 160.720 393.300 161.840 ;
  LAYER ME1 ;
  RECT 389.760 160.720 393.300 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 160.720 384.620 161.840 ;
  LAYER ME3 ;
  RECT 381.080 160.720 384.620 161.840 ;
  LAYER ME2 ;
  RECT 381.080 160.720 384.620 161.840 ;
  LAYER ME1 ;
  RECT 381.080 160.720 384.620 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 160.720 375.940 161.840 ;
  LAYER ME3 ;
  RECT 372.400 160.720 375.940 161.840 ;
  LAYER ME2 ;
  RECT 372.400 160.720 375.940 161.840 ;
  LAYER ME1 ;
  RECT 372.400 160.720 375.940 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 160.720 367.260 161.840 ;
  LAYER ME3 ;
  RECT 363.720 160.720 367.260 161.840 ;
  LAYER ME2 ;
  RECT 363.720 160.720 367.260 161.840 ;
  LAYER ME1 ;
  RECT 363.720 160.720 367.260 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 160.720 358.580 161.840 ;
  LAYER ME3 ;
  RECT 355.040 160.720 358.580 161.840 ;
  LAYER ME2 ;
  RECT 355.040 160.720 358.580 161.840 ;
  LAYER ME1 ;
  RECT 355.040 160.720 358.580 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 160.720 315.180 161.840 ;
  LAYER ME3 ;
  RECT 311.640 160.720 315.180 161.840 ;
  LAYER ME2 ;
  RECT 311.640 160.720 315.180 161.840 ;
  LAYER ME1 ;
  RECT 311.640 160.720 315.180 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 160.720 306.500 161.840 ;
  LAYER ME3 ;
  RECT 302.960 160.720 306.500 161.840 ;
  LAYER ME2 ;
  RECT 302.960 160.720 306.500 161.840 ;
  LAYER ME1 ;
  RECT 302.960 160.720 306.500 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 160.720 297.820 161.840 ;
  LAYER ME3 ;
  RECT 294.280 160.720 297.820 161.840 ;
  LAYER ME2 ;
  RECT 294.280 160.720 297.820 161.840 ;
  LAYER ME1 ;
  RECT 294.280 160.720 297.820 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 160.720 289.140 161.840 ;
  LAYER ME3 ;
  RECT 285.600 160.720 289.140 161.840 ;
  LAYER ME2 ;
  RECT 285.600 160.720 289.140 161.840 ;
  LAYER ME1 ;
  RECT 285.600 160.720 289.140 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 160.720 280.460 161.840 ;
  LAYER ME3 ;
  RECT 276.920 160.720 280.460 161.840 ;
  LAYER ME2 ;
  RECT 276.920 160.720 280.460 161.840 ;
  LAYER ME1 ;
  RECT 276.920 160.720 280.460 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 160.720 271.780 161.840 ;
  LAYER ME3 ;
  RECT 268.240 160.720 271.780 161.840 ;
  LAYER ME2 ;
  RECT 268.240 160.720 271.780 161.840 ;
  LAYER ME1 ;
  RECT 268.240 160.720 271.780 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 160.720 228.380 161.840 ;
  LAYER ME3 ;
  RECT 224.840 160.720 228.380 161.840 ;
  LAYER ME2 ;
  RECT 224.840 160.720 228.380 161.840 ;
  LAYER ME1 ;
  RECT 224.840 160.720 228.380 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 160.720 219.700 161.840 ;
  LAYER ME3 ;
  RECT 216.160 160.720 219.700 161.840 ;
  LAYER ME2 ;
  RECT 216.160 160.720 219.700 161.840 ;
  LAYER ME1 ;
  RECT 216.160 160.720 219.700 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 160.720 211.020 161.840 ;
  LAYER ME3 ;
  RECT 207.480 160.720 211.020 161.840 ;
  LAYER ME2 ;
  RECT 207.480 160.720 211.020 161.840 ;
  LAYER ME1 ;
  RECT 207.480 160.720 211.020 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 160.720 202.340 161.840 ;
  LAYER ME3 ;
  RECT 198.800 160.720 202.340 161.840 ;
  LAYER ME2 ;
  RECT 198.800 160.720 202.340 161.840 ;
  LAYER ME1 ;
  RECT 198.800 160.720 202.340 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 160.720 193.660 161.840 ;
  LAYER ME3 ;
  RECT 190.120 160.720 193.660 161.840 ;
  LAYER ME2 ;
  RECT 190.120 160.720 193.660 161.840 ;
  LAYER ME1 ;
  RECT 190.120 160.720 193.660 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 160.720 184.980 161.840 ;
  LAYER ME3 ;
  RECT 181.440 160.720 184.980 161.840 ;
  LAYER ME2 ;
  RECT 181.440 160.720 184.980 161.840 ;
  LAYER ME1 ;
  RECT 181.440 160.720 184.980 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 160.720 141.580 161.840 ;
  LAYER ME3 ;
  RECT 138.040 160.720 141.580 161.840 ;
  LAYER ME2 ;
  RECT 138.040 160.720 141.580 161.840 ;
  LAYER ME1 ;
  RECT 138.040 160.720 141.580 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 160.720 132.900 161.840 ;
  LAYER ME3 ;
  RECT 129.360 160.720 132.900 161.840 ;
  LAYER ME2 ;
  RECT 129.360 160.720 132.900 161.840 ;
  LAYER ME1 ;
  RECT 129.360 160.720 132.900 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 160.720 124.220 161.840 ;
  LAYER ME3 ;
  RECT 120.680 160.720 124.220 161.840 ;
  LAYER ME2 ;
  RECT 120.680 160.720 124.220 161.840 ;
  LAYER ME1 ;
  RECT 120.680 160.720 124.220 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 160.720 115.540 161.840 ;
  LAYER ME3 ;
  RECT 112.000 160.720 115.540 161.840 ;
  LAYER ME2 ;
  RECT 112.000 160.720 115.540 161.840 ;
  LAYER ME1 ;
  RECT 112.000 160.720 115.540 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 160.720 106.860 161.840 ;
  LAYER ME3 ;
  RECT 103.320 160.720 106.860 161.840 ;
  LAYER ME2 ;
  RECT 103.320 160.720 106.860 161.840 ;
  LAYER ME1 ;
  RECT 103.320 160.720 106.860 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 160.720 98.180 161.840 ;
  LAYER ME3 ;
  RECT 94.640 160.720 98.180 161.840 ;
  LAYER ME2 ;
  RECT 94.640 160.720 98.180 161.840 ;
  LAYER ME1 ;
  RECT 94.640 160.720 98.180 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 160.720 54.780 161.840 ;
  LAYER ME3 ;
  RECT 51.240 160.720 54.780 161.840 ;
  LAYER ME2 ;
  RECT 51.240 160.720 54.780 161.840 ;
  LAYER ME1 ;
  RECT 51.240 160.720 54.780 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 160.720 46.100 161.840 ;
  LAYER ME3 ;
  RECT 42.560 160.720 46.100 161.840 ;
  LAYER ME2 ;
  RECT 42.560 160.720 46.100 161.840 ;
  LAYER ME1 ;
  RECT 42.560 160.720 46.100 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 160.720 37.420 161.840 ;
  LAYER ME3 ;
  RECT 33.880 160.720 37.420 161.840 ;
  LAYER ME2 ;
  RECT 33.880 160.720 37.420 161.840 ;
  LAYER ME1 ;
  RECT 33.880 160.720 37.420 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 160.720 28.740 161.840 ;
  LAYER ME3 ;
  RECT 25.200 160.720 28.740 161.840 ;
  LAYER ME2 ;
  RECT 25.200 160.720 28.740 161.840 ;
  LAYER ME1 ;
  RECT 25.200 160.720 28.740 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 160.720 20.060 161.840 ;
  LAYER ME3 ;
  RECT 16.520 160.720 20.060 161.840 ;
  LAYER ME2 ;
  RECT 16.520 160.720 20.060 161.840 ;
  LAYER ME1 ;
  RECT 16.520 160.720 20.060 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 160.720 11.380 161.840 ;
  LAYER ME3 ;
  RECT 7.840 160.720 11.380 161.840 ;
  LAYER ME2 ;
  RECT 7.840 160.720 11.380 161.840 ;
  LAYER ME1 ;
  RECT 7.840 160.720 11.380 161.840 ;
 END
 PORT
  LAYER ME4 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME3 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME2 ;
  RECT 557.780 0.000 561.320 1.120 ;
  LAYER ME1 ;
  RECT 557.780 0.000 561.320 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME3 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME2 ;
  RECT 536.080 0.000 539.620 1.120 ;
  LAYER ME1 ;
  RECT 536.080 0.000 539.620 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME3 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME2 ;
  RECT 509.420 0.000 512.960 1.120 ;
  LAYER ME1 ;
  RECT 509.420 0.000 512.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME3 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME2 ;
  RECT 492.680 0.000 496.220 1.120 ;
  LAYER ME1 ;
  RECT 492.680 0.000 496.220 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME3 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME2 ;
  RECT 466.020 0.000 469.560 1.120 ;
  LAYER ME1 ;
  RECT 466.020 0.000 469.560 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME3 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME2 ;
  RECT 444.320 0.000 447.860 1.120 ;
  LAYER ME1 ;
  RECT 444.320 0.000 447.860 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER ME3 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER ME2 ;
  RECT 335.200 0.000 338.740 1.120 ;
  LAYER ME1 ;
  RECT 335.200 0.000 338.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER ME3 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER ME2 ;
  RECT 313.500 0.000 317.040 1.120 ;
  LAYER ME1 ;
  RECT 313.500 0.000 317.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 296.140 0.000 299.680 1.120 ;
  LAYER ME3 ;
  RECT 296.140 0.000 299.680 1.120 ;
  LAYER ME2 ;
  RECT 296.140 0.000 299.680 1.120 ;
  LAYER ME1 ;
  RECT 296.140 0.000 299.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME3 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME2 ;
  RECT 283.120 0.000 286.660 1.120 ;
  LAYER ME1 ;
  RECT 283.120 0.000 286.660 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME3 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME2 ;
  RECT 261.420 0.000 264.960 1.120 ;
  LAYER ME1 ;
  RECT 261.420 0.000 264.960 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME3 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME2 ;
  RECT 239.720 0.000 243.260 1.120 ;
  LAYER ME1 ;
  RECT 239.720 0.000 243.260 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO39
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME3 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME2 ;
  RECT 641.760 0.000 642.880 1.120 ;
  LAYER ME1 ;
  RECT 641.760 0.000 642.880 1.120 ;
 END
END DO39
PIN DI39
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME3 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME2 ;
  RECT 633.700 0.000 634.820 1.120 ;
  LAYER ME1 ;
  RECT 633.700 0.000 634.820 1.120 ;
 END
END DI39
PIN DO38
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME3 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME2 ;
  RECT 628.740 0.000 629.860 1.120 ;
  LAYER ME1 ;
  RECT 628.740 0.000 629.860 1.120 ;
 END
END DO38
PIN DI38
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME3 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME2 ;
  RECT 620.060 0.000 621.180 1.120 ;
  LAYER ME1 ;
  RECT 620.060 0.000 621.180 1.120 ;
 END
END DI38
PIN DO37
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME3 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME2 ;
  RECT 612.000 0.000 613.120 1.120 ;
  LAYER ME1 ;
  RECT 612.000 0.000 613.120 1.120 ;
 END
END DO37
PIN DI37
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME3 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME2 ;
  RECT 603.320 0.000 604.440 1.120 ;
  LAYER ME1 ;
  RECT 603.320 0.000 604.440 1.120 ;
 END
END DI37
PIN DO36
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME3 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME2 ;
  RECT 598.360 0.000 599.480 1.120 ;
  LAYER ME1 ;
  RECT 598.360 0.000 599.480 1.120 ;
 END
END DO36
PIN DI36
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME3 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME2 ;
  RECT 590.300 0.000 591.420 1.120 ;
  LAYER ME1 ;
  RECT 590.300 0.000 591.420 1.120 ;
 END
END DI36
PIN DO35
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME3 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME2 ;
  RECT 585.340 0.000 586.460 1.120 ;
  LAYER ME1 ;
  RECT 585.340 0.000 586.460 1.120 ;
 END
END DO35
PIN DI35
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME3 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME2 ;
  RECT 576.660 0.000 577.780 1.120 ;
  LAYER ME1 ;
  RECT 576.660 0.000 577.780 1.120 ;
 END
END DI35
PIN DO34
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME3 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME2 ;
  RECT 572.320 0.000 573.440 1.120 ;
  LAYER ME1 ;
  RECT 572.320 0.000 573.440 1.120 ;
 END
END DO34
PIN DI34
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME3 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME2 ;
  RECT 563.640 0.000 564.760 1.120 ;
  LAYER ME1 ;
  RECT 563.640 0.000 564.760 1.120 ;
 END
END DI34
PIN DO33
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME3 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME2 ;
  RECT 555.580 0.000 556.700 1.120 ;
  LAYER ME1 ;
  RECT 555.580 0.000 556.700 1.120 ;
 END
END DO33
PIN DI33
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME3 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME2 ;
  RECT 546.900 0.000 548.020 1.120 ;
  LAYER ME1 ;
  RECT 546.900 0.000 548.020 1.120 ;
 END
END DI33
PIN DO32
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME3 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME2 ;
  RECT 541.940 0.000 543.060 1.120 ;
  LAYER ME1 ;
  RECT 541.940 0.000 543.060 1.120 ;
 END
END DO32
PIN DI32
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME3 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME2 ;
  RECT 533.880 0.000 535.000 1.120 ;
  LAYER ME1 ;
  RECT 533.880 0.000 535.000 1.120 ;
 END
END DI32
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME3 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME2 ;
  RECT 528.920 0.000 530.040 1.120 ;
  LAYER ME1 ;
  RECT 528.920 0.000 530.040 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME3 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME2 ;
  RECT 520.240 0.000 521.360 1.120 ;
  LAYER ME1 ;
  RECT 520.240 0.000 521.360 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME3 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME2 ;
  RECT 515.280 0.000 516.400 1.120 ;
  LAYER ME1 ;
  RECT 515.280 0.000 516.400 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME3 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME2 ;
  RECT 507.220 0.000 508.340 1.120 ;
  LAYER ME1 ;
  RECT 507.220 0.000 508.340 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME3 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME2 ;
  RECT 498.540 0.000 499.660 1.120 ;
  LAYER ME1 ;
  RECT 498.540 0.000 499.660 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME3 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME2 ;
  RECT 490.480 0.000 491.600 1.120 ;
  LAYER ME1 ;
  RECT 490.480 0.000 491.600 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME3 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME2 ;
  RECT 485.520 0.000 486.640 1.120 ;
  LAYER ME1 ;
  RECT 485.520 0.000 486.640 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME3 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME2 ;
  RECT 477.460 0.000 478.580 1.120 ;
  LAYER ME1 ;
  RECT 477.460 0.000 478.580 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME3 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME2 ;
  RECT 472.500 0.000 473.620 1.120 ;
  LAYER ME1 ;
  RECT 472.500 0.000 473.620 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME3 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME2 ;
  RECT 463.820 0.000 464.940 1.120 ;
  LAYER ME1 ;
  RECT 463.820 0.000 464.940 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME3 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME2 ;
  RECT 458.860 0.000 459.980 1.120 ;
  LAYER ME1 ;
  RECT 458.860 0.000 459.980 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME3 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME2 ;
  RECT 450.800 0.000 451.920 1.120 ;
  LAYER ME1 ;
  RECT 450.800 0.000 451.920 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME3 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME2 ;
  RECT 442.120 0.000 443.240 1.120 ;
  LAYER ME1 ;
  RECT 442.120 0.000 443.240 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME3 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME2 ;
  RECT 434.060 0.000 435.180 1.120 ;
  LAYER ME1 ;
  RECT 434.060 0.000 435.180 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME3 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME2 ;
  RECT 429.100 0.000 430.220 1.120 ;
  LAYER ME1 ;
  RECT 429.100 0.000 430.220 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME3 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME2 ;
  RECT 420.420 0.000 421.540 1.120 ;
  LAYER ME1 ;
  RECT 420.420 0.000 421.540 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME3 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME2 ;
  RECT 415.460 0.000 416.580 1.120 ;
  LAYER ME1 ;
  RECT 415.460 0.000 416.580 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME3 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME2 ;
  RECT 407.400 0.000 408.520 1.120 ;
  LAYER ME1 ;
  RECT 407.400 0.000 408.520 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME3 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME2 ;
  RECT 402.440 0.000 403.560 1.120 ;
  LAYER ME1 ;
  RECT 402.440 0.000 403.560 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME3 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME2 ;
  RECT 394.380 0.000 395.500 1.120 ;
  LAYER ME1 ;
  RECT 394.380 0.000 395.500 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME3 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME2 ;
  RECT 385.700 0.000 386.820 1.120 ;
  LAYER ME1 ;
  RECT 385.700 0.000 386.820 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME3 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME2 ;
  RECT 377.640 0.000 378.760 1.120 ;
  LAYER ME1 ;
  RECT 377.640 0.000 378.760 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME3 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME2 ;
  RECT 372.680 0.000 373.800 1.120 ;
  LAYER ME1 ;
  RECT 372.680 0.000 373.800 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME3 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME2 ;
  RECT 364.000 0.000 365.120 1.120 ;
  LAYER ME1 ;
  RECT 364.000 0.000 365.120 1.120 ;
 END
END DI20
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 358.420 0.000 359.540 1.120 ;
  LAYER ME3 ;
  RECT 358.420 0.000 359.540 1.120 ;
  LAYER ME2 ;
  RECT 358.420 0.000 359.540 1.120 ;
  LAYER ME1 ;
  RECT 358.420 0.000 359.540 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME3 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME2 ;
  RECT 356.560 0.000 357.680 1.120 ;
  LAYER ME1 ;
  RECT 356.560 0.000 357.680 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER ME3 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER ME2 ;
  RECT 351.600 0.000 352.720 1.120 ;
  LAYER ME1 ;
  RECT 351.600 0.000 352.720 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 349.740 0.000 350.860 1.120 ;
  LAYER ME3 ;
  RECT 349.740 0.000 350.860 1.120 ;
  LAYER ME2 ;
  RECT 349.740 0.000 350.860 1.120 ;
  LAYER ME1 ;
  RECT 349.740 0.000 350.860 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER ME3 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER ME2 ;
  RECT 328.660 0.000 329.780 1.120 ;
  LAYER ME1 ;
  RECT 328.660 0.000 329.780 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 325.560 0.000 326.680 1.120 ;
  LAYER ME3 ;
  RECT 325.560 0.000 326.680 1.120 ;
  LAYER ME2 ;
  RECT 325.560 0.000 326.680 1.120 ;
  LAYER ME1 ;
  RECT 325.560 0.000 326.680 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER ME3 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER ME2 ;
  RECT 323.080 0.000 324.200 1.120 ;
  LAYER ME1 ;
  RECT 323.080 0.000 324.200 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME3 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME2 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME1 ;
  RECT 318.740 0.000 319.860 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 311.300 0.000 312.420 1.120 ;
  LAYER ME3 ;
  RECT 311.300 0.000 312.420 1.120 ;
  LAYER ME2 ;
  RECT 311.300 0.000 312.420 1.120 ;
  LAYER ME1 ;
  RECT 311.300 0.000 312.420 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME3 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME2 ;
  RECT 308.200 0.000 309.320 1.120 ;
  LAYER ME1 ;
  RECT 308.200 0.000 309.320 1.120 ;
 END
END A5
PIN A6
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER ME3 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER ME2 ;
  RECT 300.760 0.000 301.880 1.120 ;
  LAYER ME1 ;
  RECT 300.760 0.000 301.880 1.120 ;
 END
END A6
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME3 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME2 ;
  RECT 280.920 0.000 282.040 1.120 ;
  LAYER ME1 ;
  RECT 280.920 0.000 282.040 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME3 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME2 ;
  RECT 275.960 0.000 277.080 1.120 ;
  LAYER ME1 ;
  RECT 275.960 0.000 277.080 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME3 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME2 ;
  RECT 267.900 0.000 269.020 1.120 ;
  LAYER ME1 ;
  RECT 267.900 0.000 269.020 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME3 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME2 ;
  RECT 259.220 0.000 260.340 1.120 ;
  LAYER ME1 ;
  RECT 259.220 0.000 260.340 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME3 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME2 ;
  RECT 251.160 0.000 252.280 1.120 ;
  LAYER ME1 ;
  RECT 251.160 0.000 252.280 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME3 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME2 ;
  RECT 246.200 0.000 247.320 1.120 ;
  LAYER ME1 ;
  RECT 246.200 0.000 247.320 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME3 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME2 ;
  RECT 237.520 0.000 238.640 1.120 ;
  LAYER ME1 ;
  RECT 237.520 0.000 238.640 1.120 ;
 END
END DI16
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER VI1 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER VI2 ;
  RECT 0.000 0.140 655.340 161.840 ;
  LAYER VI3 ;
  RECT 0.000 0.140 655.340 161.840 ;
END
END mem_ker
END LIBRARY



