`define CYCLE_TIME 45.0

module PATTERN
`protected
U=42aVVbP;b[gHN<OKZ.;ARAKfYEMX990\LI[[0dATB1A&A&YFBK,)KM#T.>5ZF(
af\,XGO:XPW(]eBf/Q+7I.NF3,M2L55gRU61+/RZ9GY&OCK^+(M=WUIfL56L/BR?
M.V]bHUAQRB]DS7Ke7L>C[>V@3V(9[M1eNE,AY]3f4F5aA7]JG0SX5=519XMfKX?
b=V-1B2<^;,Lg\YL+D?AT;XQ9:O74_.7(]EEIX-Q&IJRD:/&9&R/J&>N6E@(He)/
b.[eD_(8//S]He/T+S7&QAIGK@B.?g+T?DK:4Y:-2O.CF78<2)7aH61]GOZ3GJ#G
Je/f@K&\3R?E,F4NNP\b^/(,UQZSA6J1L^8TFK962G_)5,RdU3e,fLAZ]9>a8&\U
g@:7&/13=geZ?A/@[T</S/>KD.4ed6f_d#FAR:JDfYNUBc<d9KJJ9G5_2][DD9O7
L1c]:cB.QGK(#KHLA/PSY0c0c:V5S/&[X:\GCaa/#PfTYJI@DZB=d)8fG3[>[#GA
c6HI8DYf_E[STR?JZDa+5[-XPZ7&99W4]aB]Aea3g0QA3CH9]d6R@?0fDN4KZ.,Q
C1Rc8^@CJTXPH;F9>R2\g.(74_DP>2?]W(7Z\\GDXGV5MJc,#=9J81>.2C@?2VDL
[#\8d//)a,Y4?O^6<A#c]HI6)QaPU@R-4BA.N\5#OCPGY_\TAK<H[9/L+#7,@0L\
(3XG0Z&P@@^)P+R+=W6I?(7VT[+HIM+&,9E^gK3b9?b3N8##L-(&[@R.8DO]dF-\
TM@K=OTJ:F9H>=&_a,N<4WBGBT:baacRH9O9P22;MME(9aR_DSS0<5W2_QD^f<P3
7HCPPC23HG)/+WL[VYYL[>XD8FcV-5d/J-;?NU]H3((;9\[1^)^=@WQf8FY>[d.R
Mda;L?-R,JO?4;bO-]ET(<6_K4aa,Y75G2R93]4YPTHfTIF==N_(Aa4bN8O<R35H
3D.A(O.9H/-[<+T-KgGMB?#dXO>&7DMILF]5760&5-B&.D&BST9UC]&2Y[@(_H,0
9Sb7-Df]eX^G9:SHE6TTY7J2X-(N@NK>6\[F64-+OM\2M0<]NF:U6V:#?N54V(9T
L[[]YaAL5fBGXfS<f1@H:DS<@E#18-b1T?[3.?,W#6=-H@P4Y6dIK(C+N]Q7.[]3
9DI4WHLA,WEX&JA?V(Q5c_Y:UN3g1=@AN<E]/+g.QZb]c/DK2<,K(94cZ)ZSL23^
HQI=K\IOdR1bF?[QXU2(8MB77c1_GU&7U?N#WY@E8G?U004G@_K1V^b_&A?7UET6
G.;af/R?+D8U+^Z+fG_S_=9gKDOOaR:?+Q>QY0:-\LPW-.7&b;eGJB5/0>ef2W0H
9KeZfVKYKV/OT.f3=3a5=L^YG:6O6V.EW)6#>e.@T6R0>fIPgBV^TMVEfD.gNdgU
^-75Sd/@g_;JNA64FW\X,JAf;b^8XT69(9C#e=BF^.&]5?2W57-5S8(0WXLgd_X7
M3Z?F4.X<E7X2Z4)Ac;;GV<:0gA9=12TKUTJUB:Q+QNBR.PMO<T/FOP&V6,;5TA7
XVb7CU6[?77DC+5<6]@]4[9M(Ff+#(JJce2QZX&D7Q/X@5C&<f]NU]??R\=E+E=f
)N?4B]fS,3f#]<WDRbUf4^\4-]2V+4E,UU.CV)SYDZNV\\e,5=U8WYALZLYD=,K_
+6aL3RVU@8QeDMA.XJD1ag6YL[QOQ@bCadN2C5T_JW?Z+K-U@=-DY),P+_1Og7:.
VZ2K;&V[JCBgX0I>U?#TUAA##G9EE[62NWLBW?SK1e+.A?.V78X[F9.SJ69cS(HH
,?[Ag)f(AFCASX?YXBXL6+6MMd62<dTdN<BINWC&:D8Z7J+Y-^5g066B;0D5Xg_N
0V)J=U]7M9^Ud(>GQCdSB1;P,Ad:EED<ef#?)a31K:)#M5>,(,HQX,XO:ZCBB>&1
eT-ZMYRT;/K0L?8E0]NbUZ[3PADON.3GYJ_C&/I/(e._ZZV[Fa;Y/:U,#\\4[-\9
VS\;a+g5SQM1NAa0CAKBRePf^LXgAgO/-]Zab]5cd=MKC9\8]B7A,E=(7X<UHa7A
5I[,dW>UPXPaZPAPAO;F52g#X(Ng,2>e&1S0SCTN8A70BJNAZ.d=08=G)K#:>#<_
0Z7^X38FITWKfZNQ]H+.>LO2K(a1.I&aIKS6dZWMQVeUK201)><;aQ):I+0QOC8Y
^FgU+L>J9V:.,HF/2C?)3d7#b6)RB@000ffFITU/J7=dW]T(=^61fC;-.?Q]=1?@
gBf]\C2UV&.fQ:AH#G;TJ[PX0)PWWC\\@@OK4S2JAH6)-O5XB?PF:>eZEX124^ZF
_EQ/cGgPYDGFFU5E=^\SX+>I;0A2PR_=J84a7cQg(VgB+fbBN>&VX_-Xd;R=ZLRU
&^5LU?E[FE5=d5/McRX^Ba4F[VV0)663JYC(YV@;E2Q0dOKY?23FFKbc4U73Be[C
2((2eVS84;DAb@EH0E<b1,HHE&7RfUcHKBC/5^/e>[W#OZZN5#VffU\Z?4DfMbC\
I<LWJ=76_RZF#JP6Y[P(0bgD_Y_^-HW?W,:#2MK?7N+T_<LO:=N04<9AL512Q8TD
U;b@RF];IDD9>2_,#cARL;,a1RNR/#/OUP:;(/F1,N).L#Tg_?a:N:V5O:LH2#C_
9TQVB=HQ1D\LY0X#GEM])ceHe>[MId4N3:?V2cZdO<8#M9[RS-OKZ>XK]&I5LB>Q
@.D)c:[984UP>&ZH@))YQ]:G\W;B9@ROY_U,HWU09eJSdX\73AXaeR<GgZKd71,7
?DM)E\.dYD9W:E+;28I#73#S:37Lb145c8]S_J=&=XXB>U(Qe(3GG71LL6F1FE]Q
F#WZU<(UP8If0TNd_HH,>:[:FYEgK(T,b1e_/fL6EN4aXb4<F8W^bA5F5P)KWaOX
+Z7D_GL202d2Ja-5AaZ+J=G^<=2^d=,0Z4X^1CUAe0M2c+6fG?1O9)-[0/(YS+3_
Ua:ZRT0M@]V5O;3N]_2TU4=IMEcc>P]AI]SN1)_1;?)IDBIXcL-?=]KJddIX2LVC
6V0)>33U[53Y2/N@+eZ6e>3aFG_1Xb+34YH4KS/b3WI3W1UL=Z)F,WfAD<FTY(NR
@SVU57:&I9:TNC=SEW34;<U@eGQ3D/&BT1@IQ3e@::aB/e&\EY]H5N4K_3.N)Y(Z
O8:-eCYe/\=/AMMa@LNX\1-<02<e&?JUL\U.K4c8Qbd(Y.GU.1aWeK39F-I;aX,H
<:G7VB;B\/6EcVc_^&S8bL_ME0#L?64@GZE_L)>TQVSN9#I#Z;Rb3e0fE/.KB37Z
d4CUV4Zf<?/Ye[AONL8^/.Z/U1XX51?#(<FRE_8K#g3PG.&VHQ>_XZK2d[(Pg_>9
)f[<Ya[bBLW?0E<T.MS>BLf)fZY_Y739^<13c;c2P>C]UaEXY.W.?:C]7P-]f9+-
d.>B,FC8LR&DB3-B6Y2<7#=KYe;NUWDFS::a8FLf,aa+(G##,8(;;:J+6IZ5Od71
d1,^=-PN-[3[[eV2A2O,KJZ]d:Y.@.Y^#bN(?7RV?M;cP]I]AAQ@gaV]/Ne[6XVN
:PWcW45B#4.M8ME?RPT:d:6&7PE4;/V]::b=ge5J+cFZNO;=Fe=L@<b4U8K]bc3<
^T^g9V0\^_1>ZWH@f.;OHU9fSe0@)/dS[?<LF,V#(C\.A/9&DcZ\.7+@E;JV&M;L
bbf.Z:a[][7B8G:aETCGV.ECU/Gc&.M5gIK.D]YfN/d3]C/8#+_2&S/<I(>[L#/N
DERQ=XV?^>(26#T35KXQg+XBEUU:<H46Ha1U@)3ffFTTU6C5e1IFVQ[R6A3BZESP
M)8KH5>PMGF863K##,22LT;5R9[_80V32V(E#E=<H=#XK3ZS:#V;Dc,,<Lfae_[R
8A&fYN6_JOFY:MYPU>GKe?R-7D02bQ08UJH[(HeTVY^LZ+RVMY<:)^X:Ig](D[JV
@,F[&QgCB^I27&Z<B94TO8XN4@59-8+8Sd&1eX_2F=U:eDB^BT\0&PL32CI?d84L
8?;#g2FceI][&JQcNIdgHM3SUZK:/J4^?U?51D)1#Jd61eI0)H55Ec/3Lb=)gg/+
OEAJS/B8KT3d-Y8I<.^2X=)b3[,B7]5)b[?0_,5/3OTYD#6DgTKOgd=<OB=P/#MG
A,^]KSWO#5N.GS1M3838RaFC.O#X?)4B7(NcF@+d7+?TD)(3/22(152aSQ+/I1E8
)1g3.QX-XcOT+L??U5.Z?W8-;_\Od4bBZ_Xa:VVHXJ2]@P4Z1(,2[(.#\4NS/=@D
dUM#][9RUFA#XFg^:;b?>B/1(gEN.Z12F&<bIXY_O46<&(9eRRVK<KMMF0@+FN<&
?;O9KPW9XMRc3O_7[+A-P)0F>Y5.76<.]6^?F_,/O&?bgQU&?J67VcA<1PW:-(24
5;QWg0NWN_V&:&KNAgL;6EgG&01M=fN^_7,9^@L1CRW)YC7K@VVAdgG5Q<YEC?ef
aPVU]<cSe<CXf.?4#/GZ(V=/[#eJd#VU1#NYTI-^@)dXSC:Y/XDHg@FYf]2V-Ta#
1XNU3>(WE^aH#c,d9U#g#4.X6f9X+58594+>8C:/[XPa0>XWL9YOZ<;A@d/>3YBG
W3YV--fC]?>PI3(R79V/4RC2UM@H-c[:@F--S^Q#AMB0EK.@bR6&F+^>.-0;B41[
8^MN</[aS(IQa>B[#<c:G_68Ba)dVeGUO23B_<2+Kb>0D4M?:ZbUbF5H(5[?W(O:
J+?JS_-^IT?1f[gcNSO/MWR>M@eWLK>D+P5/5dDfAFQOUG_2H?=?/3T0C#@<]-ER
OfH6DAY4H0SK3_/0(XfEX4[-.cJc.R-]3]U)(IPMD=fUI19PY@EP(D@NL9P=&4@^
DN&I1;:MC1]6I.MESePc]OWOUdHA^EeF4UNEbSc-&VDH^/JDU0DQ/4=J7[g2&#+Q
LXb]+ZL.16TR^UT8&A^1Q216^Ig=_^+g><<]P4&GL-W+5.5ea3H#;O^80F(?DW?)
AKTT[c.ZT&8I6UD,M/):/+Y8(P^-?O</TB&9MLE.5e?c0e)B5A.b](;HUG/-4Ae<
]aHd(:YL)5M#_H\D\VDOPBJK>KH(^#BO6=DEgBY]#.+8A(\@b3:5[.LgIWU\L6SU
9<CeXf?bW6\GNDaP?WeQ/D3/(2HF(:L]C&>;/P7gW>Ib5,XZPDR?=34QU5g^#a/4
MZd]2T(I/U0(_8^[M)9=+5?SGZH]>15V6:;9KNX97#>&(>X]Md+<&9M/2b8MMN&G
@,+S73J:,B7QM/M6S/5.V?&WL9V4H.BfHfHT8AJ4a_Qa.Ea6QXGf]XCJ[0>(2=J2
7b-fN4R4/:9Y,JDJ6<XZf2BKSWbS=7,PeS/WfJF4(@c3JN:+CEbRQWc;;:C6ZXA>
T.I_60]eQaO.Df1IS;3/=Y;GW0U<A;9Z_+8K>5&C-3cH76@71FB=Bg(:Z)8CBY)T
bST<DZb=cKM,[H(^E\9^RbA/dO<_4UQGO3)AP;9S]PR.+<35N)RPL(/URYOZDNXI
M)1A00b:FV;9UI#(@MUJ/M4/>;4<QY)KUTOc[L0Ta)X:MG\N1A[?M8,HI:N4_6bA
K]<CZE=^[fG=#=4HUaeJN:8c&>0^:4J-QH:YFE(HBf[dfOQLH<#)@&;F;VOIa(<4
c@+D^KN19PXQ72C=L;3gJDX8cZGNZVH+7GM6&<[cOfP#cDbD>5-RY@&=+U@&+e+_
cHc0)S[STS?S;V/+B<b>-/GM87eLa2/Q_:]8XgN0[H2P<C7D8E?#]\?3(6ERb\9=
VbW;RYQ<W9/HDT38;Z=f3[cR?M44TP4;+&.XH;RYOb/,VLHcNDG0][\W7Y<RPb>V
Y#H>:#4G>,TE+eUY-XZJ8;f8:KY(=5WPa=Ne:4gI.]Nd]VHAGaNYTIEGfE1,.K=J
4<@c[(#+8NO9C@9))Z1+5AR1<Ua_\(/&IS<6gNX#1>\J0,A9)I/O(9d2J59>[U/#
Y,R@I8(eGDbCUY^/]OeG;[VE#bXa20Zg2?=(HfC@Na&R;e-bV1Z(#SW41dLIRYQY
3@WT)PX:L6[ZeT7BQTDK?E#^S0aQGG/;^E=J5]bGNRcM9XC,bAbKEC/9K\@=Iec3
DHCZ.HGVXI.\\RLa-&(A:K@^]9.NM<gJcGc37J]c;B(-+V7QUS94.4;1J@]_-OSa
9=3HR.&Y2[2AEJFLD.D^Yd@F3L9.C2#bfFL12>-_4SJI@<-(>WfY8W<<_12UF,Q)
aP6,d@)N2G>S(3A[NP+E-LOV7&XC7_,9F\<(]cd(KL3R[7BHK/K\/ab\\EMOa:[<
GWEAT<NBBTA&;+eDPfI</?QR@2[9IgTg9L>-BO-)@<=dO[,R5d2MQJ<Z];JaGUZ9
0/WL,b5N1HcU1aKb#;.<fRQ1_(XfDa6@[DQQe[dU[=Y.;6WBcMUTA:VO3<LRV<W<
=ZNeL-W.C?N2^^:F?&]N;IHVTAZ06:U@g1VfB>OG#ZU1W3[-=5RA;>bY9f8PO\^M
09U;Ef17b6\72FY##=^PBDO9]cGXWcaEO;^bWJY7OFMf]2HIV.(J.[#bD6^?[PRK
b_;)8^LA6=FbBXf</Y#d<:@Ga=cdML;=AR(1#U7U-(>9/DW9@YM48M(W\.bF^;D#
LHdBV_YJV:W]J/HQ>P+fdU)8+FJ>?eCaB[(IVM9U]E_4_P&;/Sf@:F8M4,C8A/GM
Ge8ceE[LEGJ2^ZX:g70<HD^(#/X^[cf0_aAaKAQa<A7=W?W6AND^5B.WW,OPBO5H
,L:/8g)FZHM5M_-Z1c1P/a>7MR<26FdILIQKPTb_.Yg5_E<,C?+JD0W#02f0=4H[
/b&NW?X;<.Qd0&<[B\37;cO/N:\cc6Je]YdS[_D)+[:2^(.)>bFAZXO.2?L1C.J&
HO^BCP3F@N@Xc=0A)#/J[)95<T2Fd<(H+WS.8aPKOM<RPC)[EWZTTL-]f8D0_@2<
H)OJJX<IT.NQa0\47#Q5QHCLHCTMJe;6[6Ef)Ne)g<=^]^Z:JG/.(OgV+P8ULY66
#\Yd=4R8;I@a.B6X7,=D\Q(&>?AP]f;F(?X,?-OP\=0TPL0Y1\7L=T<)WCFY@;]Y
98a]X<D6bNGGG8XM\=)MCa/\&=F-ZfS5HZ#X\5]fG)UJfZ:+OER/:WF<aL3IU@P_
QHPVeCc&X)^XGKK78=G>T4.[YXM?I#P]\aZX?YT++DR[Z/a?,.U?HA=.F<#dAAOJ
@&ZRgUG^@0Ag1B8KIgF<bDJ7G0S=Y7&<J^Z16\RVBJR#1RS;+9MfbV>Wc6[6RY/)
@]0?BJa)K\e&56,E129f<LL\K;=T14U3^^UXEO,HA>@Z6f[Ia/^V0P6+UT=5)R)6
H@]:?Q,W/>)V9Q5Y16&.[8F8=A]P8#D?Y0FS+(Q3X6V4Ha&:J72;/>.0@CeZ;THD
?.##T8R=+.&?M08G2E.V;U;(\c[;R?a-V(>.KdP;QC&<S.9J=FH:SSZ(2O+Q/;X7
6;g^PR-.<8+UA]1cI^(a&aIU\HETg^Y1[V-?BU#_OH;Y\WIBS-Fa_G)G.?WR#]TU
H4Ff6+P5b[YNa>ZU[1MOc[NOJG/<6@JH(-T9f/J/3V7QLA8,(I1PKD#ZX5V(.aJ)
1.:JOZ7M<@,f-aRUbd5#L:7)]&\]@FTL4Z=Q<:AaJa<3P&98_8==1fBSZJeDPLDG
->(.XHG6P))P]5[R#DDGda.EY\G<6=fWGSMe0/c?=G3gbJKB;YE&9bQRWK2/B92N
gWd<68L3::2?<KQMY[R2NS^B1^A_?=ODSUT\bRI#g2c5K8AIX9PaFIXUQ3AY;4dX
=f[(+:Z=ab4;#gNS<W2N&aLR+8SH]d<6=G^L//FYT^V//;K1MNKb27_8[@2</G32
X-@M0WdcAM6?S7Qf;Oe6T&-A;b=e2IRFH5-=R@G.OVHBb.4<9M>I&WX2>ZW1XX)0
aP\cN^;5TfcBD8;-5f(b-2(0AXT]c)75W2W?<6ag2-b=cHYE25&,VaXe6T6CLdb=
H5W86IKX:LRR;aKfUfIV&-\MScDSf3TB\EAdM4W7c2.f#6[)V3UZKCaS9983RgdO
S<K(a<:cc20YQ03SGfG.;RF163?S+.\0AC(.W09VN@?JL)bIPSBG(2^U:@HZS/#B
OQc/#]b70+SO4J&L:C44V9U=IXD]@XRO>=9>f1<YQKY>3SZD1b\3\[8&KT48_3b:
:,R19,TMd<N4>(LB7K1P0<R_b0I<_I-9fGTHHAdbe;9I^@=+@/GF9_0@=]d^)STB
304.ga\R.SW^#f_4gKJF<;/=;L956I5EXfZ+HBQ,Q4QdT_K>2K\KVONC(He(;38Z
K&_LX9A,PQ):6c]?BHZ\VfAIV-ObL..4W/dB2Tc^Z[dQ96Lc3FP5L]9>.a@fJIWW
4?C<S=-4AI?)F2OC.G#YGLf(WB=4_HZf_@c+\@e7H=a(.D8D69(F5:Z;;&\M^2SL
W<;AXG]=\5CFD1^<HK.WDJD?GJF@-TH8[d)<2F][5X47;E&<5a1V/Dc@7ZG:C)_&
2,AO/_5d3;eF]^3>#?BG>Q&S\YgDKUFY,(9:@=(1Nf,M4eE+SG6cUN&+)XCDcL-R
4F;\Ae)OeXWd\>^4SGLF2Y\^cGJdZ[5=;P)(+L(AWIVe<&2L:VYd;EL+DYA/cO@+
ZREZ@Uc[Y-8?071G\W^2TH-1.MVF4Md7#b8U#0T5eF\I><?CR1-ZVA^;O?,F;Z;9
05Q45[CT@TbJaKUCb>\^0[A]#/>afEOf++BbRYcK/g[48A(Y&e/E1_^0-aGN@D(]
#8K)89[^<K0CBdP#dTb_QF-M+geX;KX0J:+eX^(BdC?;4=.;05)XIWT)=LZI_TBX
Z#9S-TL5\O\SLf^H<B.@)Og8AG-K+4=E7.6NaQ-#E+WF>\0Z5F9bTE7L/\\9V8D=
a,VSHC&ON(O2DF+CWOYRVEBCe4,D3A@YQ/\KVLT/#-5GVLd[XL\YSe[/;[&B@Z1;
57JC(?,Y&61-]>SP9)g#QC7XTDVOeC0:5;W-)+\a,&.eI@V_P6\]?)-bec\T8<@W
3LQB1QN7V:54Cd#6a-]fXW77R+;-Ua,S:FM_eDTce5e=/E):8J_5N7VLOeL,5PeZ
&UWX:3R]F)aUXN)+5V1E2D]b->>#MPY6EH_=AfLf)&77&<TgPI&a\Q-)-EWF>D(A
+/7D;ab2VcND<f-]RDU#.QNI7\L^@HU))M23\_P@-5N/HY(GV&F&(FN0F.R.FG8R
>G=MIXeB6=/Cf^/EXJOI)\/F+ZK-V5<+,\^6#GMD(4O?dMNZU;-AOA>V[R?0a8==
X7[+5WR,U23)7ZS33c-7.>Z]1TJTG#eTJ,-a?A;+>A=:Z/#=VgcWT@(:4&FKKc\^
&=O_BUJd[/JYeUbWdLZLD.@VYO&7F]cT\?bF@b3M,LeKaXM.G5YN5?L^IB,5-S4E
C0/Dd90;W+-I#<E.9#^\g>\d0&;H,HN<T+R9QX<[^GDGNH^@IJ:dLSS3=^M))@\@
0LIQP+BL6TY((c+2.<MAcC?&6(/@#WM<88^=NZ<>.B79Lg<U_T]U4Ge62381dd7W
9e>Y0,L8c,]ZJ(&ERg,AGHJSOD@6]6VO0Z)A)KAK,K>SG?N?-C?6N1\5[/B\X4/(
LdFb7\G1SB_F#NX4/C,R[FC,S<A?MNV,WRabWWW_2)>aUgRBVG>PY1^7B8<?VA]2
/JKX\P#?(4(HF<#?GA.?b/HR=Z\]SVQ/^WV.Fb2)[06D77:40MRECN.Z[b)(Y\\R
0,7^bA_aD]TL>1))92INL).Z4c6P>?Zf>F0,31J,W^ae#F51+6F3URP.=-P\#(8<
^.O/@9e^QXP3O@+SYWC6N2bJd[&6,ZA8e5TL?5X/E]E-M.RBNG:=;47WEJW8AgBF
]O#.UG>2MUUJ\)=3.E-+bRD7[e^DZ=H6]&X=0bBS2,R?)fVg0FfHX?7;VO6Cedb2
&d8G49&@/]W<IM]O@WL)K\&\,3IGU1G0,NgAMM>A9cCD6P\T]919e\1NC&/T&AB1
/POEXW_F;W_09?d+C=/+9bOb5eAA7@eP\;Q]gHINK1POX8(3;b4V@5^)0[Ua49WU
@R^+&WdNB(]/g?P/fZN&;U/>7>V4Og_Pa]3A?L25TU#48>PeGC\d0-Cf5ZU7HH5>
&&(;X@3RAaa&#KUUg?2>+WCfL3U0E=CfED.3@D@&=fe&TeBg?@[_:YWeA\FJ^>MP
]gXc#=[5fKX2.2#gKPA@#VdVF:@>MQSX+aff_XO:G-Ob1>Xd&fP(7.>N?-OR-f2N
aH&_8./A(7P(Zg3DQP5@e6eb4<V?.CV/5YFb_^.:^9V\PLO04g9Z[#B:_0QN,1QC
R4b5-GaI3d8)(+)<caCcQ_T9a5WJ[\^.Zg\EL+]7C^(X_^=V0aAY(gWgXe3O^fTP
],FQB\:.R:Z1158)JAHQP>7F:>[PL-CfaBEabX,.6<BU8&XAR=T8;[MeQ3=ZELLR
@Q0,dGJdE1eD?;+/R[NRcY8WW\D#R&LLDYF<_Y36)&,+:d1S1]a7P^-X#,1ZRL48
g.?Y:#BdC.a_J#fD_4dU:3[O=/f<[[;E>J^Nf;/Ma&.ZgWVLBd6Of;dP)e#/T/^8
7GYa&17OTLOeAP=08=@YLeLP#GZf79c(.7X@?2NF)HN]N43e4_[f-b2)I=H<BG0N
g9,H+058GfPD,:OU@B9LfWVTR_=]83Nd&?==1<I1)R:9?ADa6DUOSV>1_H,ETgC;
Z=gcR_1+Hc&3,Z:R:/U]SMf3GPd3Ya0Ba4.ZP7?7Ybe(IUT<:+-UF5O[.1;,3Ged
I<E<2,DP#<A7S6@L[8@(YeGV^C_M]]RSCS\IN:M@c?6Y\P@Z#R3TW@_Q3?(B.DcK
(^&<DTK04<A7&9-OSEb,c^\I/<)a#)[?g;-1^61^4aCQDR\IKAY),\1:X1E&^XU3
1A\PMW#285E;PFH4CJf.X6N=K7JG5H<P]a/KC9>4W:g=NC4ITL,FI1fW_0&:-S-a
)1NTfffR>^9.<M=KgbP6_4KOVSHJ8@V@C;O=(Y]:f5W_a9a,,:(<:CV.J7Z3P1L0
PNWO-VYYB=]_]OS]7\R_GBEUE(7W2U^dTAE/EJ;UX?+[NdS[^Q>/ZgbW1UYJ0PE-
#Q03L7dSTPB9:FEc8a3.JVMS59AG<AZ4cf=9g4.O?CRPgCT(-a]&<9WWCL->cF5V
IF;3fT?b^))YIb^/=Y+[MZBO@B2caN8V;S0\gV^.BcD9ZMfX:c?@,L:U)8QQQ9;2
Y+.FCC0=NK&ZOR0(N51SR62R/=,MgB1.0Q(QK;)+=a;.9G8#_MM_^G<0Z/d7-Y.@
EWNK^VJ<O/AD#WX)=XJ4A[eI(Kc>RD\@)DHb/bW78fH8/NOLf7QC#dJ[+,V;0_Zb
32=6-3\2N.0AfeM[;LUcC\<JP.5RW]H;-e=OB2,6ZJ5U<Y#OXC-4QWX:+<,PVG.0
D?UZY://IfL:5\Q/-:/6fESU3DB4&-FDD<+G)8SB]a<TPX^.&,0ER63/(Q^NM-B<
=?<(eN@_[gM<NGE6,&9&O[8[V])DK;JO^]6/gY#DNP0IU&Ce[71>Q<YZ@YQ#fa-S
.5ZB=SEJBQ2XX\CX&Y).+7O_?MbMGCP3B<D&cS4^]Mg)&C^bg(PAX:d3S_Ccd.W8
-=15=@]CQa:+,;Ca)I(Sa?/5;1@\bQO8J^W(=B85G@4JA+aQR,[D#/V9[Ya^)aKI
3^1OZf[K2V9RYEI,-J([BBYV7;BB-/I)C;)6:&UHfgS6_EOa4>B_#JQWEEWF9++,
W)6Z<1;(8.]<KV#&e#XNGb^FMB]G<1UfYfN984NH<LB:]J#&T6Sg.I0>T_+KT0>C
GKBMP5GY;,g<#R+:bS+8XE8^IUeP4CZ<TM+/P(A:919SYTX_)IX-?9OR#=C(DXBU
6&L.c[-9D]GTM6._EZ)Tc(B4OD0-+PRA6WS>;[MfQJV0T/OK]3&KX.YUMIbg3:6C
Z/(SLW&;(:3b3J^VfQF9cBIOB=.DFHRP4X\(c05\\<=G4BY_0JJ018V=OZ;_G-W3
31_85[H19Qa]0)GO>5=4MYeYR]&<A-DebT/YAg<E.Q;&bgWI>gMcMJ?7G5f&_\^=
ZJRCD<eQ^JIUHZ)LFC+D5SZFe+/?;.B)^af\#4e=F^U_L8@XP4(VD3)EHTfGFg^5
-3Kd)77F)JGeV\Oc/2=H4[SX?R,TZB4HW?Q,e8;c?5fUI93d\8Ae+N6#O?a/+6+J
Q&GdNPFdEfa)^=Y&a<,>MPKKR5KcZ:S\Y3&9[fC:OKM@\E_=Q82FBET15FWd:)[R
STJK1YR<ePcV?O]]CZaJS1]ZCZbXdC:XDYZ>1ZQD2&<g8cf:g6>fQ@0B5:YT-S]G
d_g6Z&(HWe1cNBObg6@,UW]4aE-cD62_560(6\f\P=(&PD,Q2#)PG.48L5#MSf_7
/.2AA552HJ7\TL9bG@a0U1^Ac]b34]WUO/6>I&[4NE-CLSZ9]d^^&_..Z9aL#efZ
c3]7P[GTK^c7R)BWeY/W]Z03B0Y@Fb1@Cd6]D8/4D15K]6=-3]ZdTY(ddIBBd=_5
=d;5[62/]Y86dM0RGTD@_^^@]e.2Kg;V61KYHc_.Y.8LfeN-.C8e/Y+S@O);fgP5
LAG?HM,Zd6:5=3Y,M_Z#.[4aA\</=9E:D6SC]73N-/Mc6IJ&T0&?gg0FQO(=NM]L
>AJ?J.Rc[9\E5,5LPca+d9DRQ_IPD[2<67W_V1XK@.X9[E1]JS43\PI@1c_g=:4R
R:YU#2Re\<::V&^Jd6T5LbbL@6\A&N6_K&FOc?Xa(ZR[e6#?)A-G4DDL4<\@Cfb:
T<dM)0:1]T=2,\^_G?fQZI?OELTU_)+\eE4N?<@0KL)V9#:A[>3W2XHA[1-8<1N3
]F/^@A.&MGAP6T330B?()?90AJDNO+70f6cBF_FA-[H1<\Oa9-Pabed-Gf8KOW2<
M61SXaS5eZ&Tc/F1\2-RfSF@I>C2CHXcTGDb[6KL@]V7=^(ZdSN@&-X/NCQ==N-U
Yc.EK:(4b:fa<3(2U46T?]HHgY_A,a)ga.4A[6U=NHFaC-fb93AIGRBA18RCH)=/
)6RN:X:Ng(X+CZfK?=4WOT5;.DCX&@OO?8OU?@>N\NZH1,RQV+@gc?P+P().+cUC
Se2M9#]_ZWF3\QgXEX-L6^-)bBX46RYe\?Z6+@M4MB2eA(f8K:P&>7#C9#TK;f<W
KMZYKeCKE.QGLdJAVU[+_GV@Lbc9JBH2][L7Xe]P/MKUCU7[ceM66fGX[>-Q/@S-
[Z^508RaAWGeOQF.QdU&4A<870M4<LY>g,=\I4ML7VMJ7.a+Hg(QA,I]&gE99e>a
V_+^aYf&9@DP/9?F<cN85@=[If?5,(b=QEME-1-e4M8\7=ZWMC#O,U3G\CV+8G=@
<4RW<R:);3=M=L;cU\>PA\aZK4R,1<8b9FD#fND7O_eWAH2W;-1QfQ<4MX&U3G8>
?&Q2?X#2)3HMGXG=^QWcKRaHTK8#KT/AEaF8/D2^&.Q4-^CFW#PS8SDC^WR<c7;O
ETfZX^C3(..C<@0+b5_VBZUN;#7H?3c;7\=DgSaU;U:30f=cS_L[I()1[CJgJTAc
0dDS7M<9@\gW3#2F:HD8d74Y^V7bF7Q^,9:POG]#-R^R]EIdAZ26;&O/g_L5A9TM
_Sg.^=^;I^fQ=g1/@;/?]CVXYD@2[3?T#-6]=T^96,(b+b:1H+XPNYe5L@UONL=<
eb.Yb@D6FgRWY@.)0Z7?T[@VO^Y7N;:BX8RVaCZ\(E=G,&&]WA2>]6>NgYgJ@RPQ
JY6a\TF]DO(.YRBa,3ATV/PP<]#Y@gA#11<[C?)\aHWE;>6QcHTfgdF=:RdVJR^=
^^dT0:5&c#.IPI/3(gDOU@R<&XPRTAg+:[cX)AaAbV&gEZf@Y9.@M]2B<a+Y9HFM
=cR^U9gf97a67(BaO7c?547@7O)MI6\/C998+J6d+X]=<.A+V8B_&DB_DWf<F)-A
<bQW\;FB&cZ8Z6&>,NA]-A/T]E]_Q:3^gU:-J4>g<CU&=SXRFTZ#HUS.KbFUR9bH
S6MI5^M7WH[H?S<PP/XS4??2B?fW\1HQ,e_1MfTOZM82f9[E0[[^Gb4g;;HCFFQ&
L/Id79SF4OTPQ>(?[6AIN&;bbB5ADNd7W7))fNE,c(8(1XeO#IL/W4UL&6,QEP=g
Rg7CX]c(??e:LOD80IDCa32XRN2+R-E0b>dI^ED3#J\eL_dXa,3Q8:bG#,\V+4/G
fV@+fFSba5W.@ad].Yf:#A.5#J;e(T-_QQWX2\Ee0(_7a;6ffX&?dF><M6Y?AG(-
6f[_-^Eec&0ZL(L[G2?Eb_0K;J4RGHa>>PTf2K7Z>EOF>)X_O[[G-<.31V7FcYbC
A)U8UMb2ad>aNgO<=E5I^HT7,c-N=8ZS/F+>[@#WfccH]>g3AOf#:A#N/\WGA,FU
)^+._bX1D38-W@0=?e@NJPL()6?47_/=M+JUR97V0GB?W1g;1C6>ZZ.YAAe3YK;c
Y:g5A4EKd\G).T5I?a3VfULX6P-=U-&(]P58(OD7D6aC8\CaETT(c&<F(C=-c]3D
:5343N3.1:KNG9#NE7\3a8gYaZP#DE?E&R[&:-ZEAeCYG<1V:]US<2@JKU]#?75R
=B_J3(Pf(3ca)>I4GWfeQ6RPR+ZSa4]3A=5^YRTXd9>ag/bQCgR6F_TO,[KD49\G
XbLf.[N(4_BM,53Y(<_9Zd)4NE4A_U;&+676&aB?G&A5;KH6\2-c9MfbLR43a.Me
b?<?&VO)=2b4Z3Y^]TdMW5/(?W#EB28Tc]Y-KGEATBR^09EPf=&[@@6:AP@+D+]D
F-1MIKbA1gC<Q@_=:?2KSY82gZ47Sf>PJ@J<eQba0aXgPIc5FT_=/>cO8505.B=5
Q0RKM.eN[IPHg>-F+@g7-MX60<S-,5);7A2H7U2@#LPYE>=]eJJ28F_aZ/J>aI5S
A6:&ELNXUJIMWZ/7YEJ(D>]FVBX:M>dB<-T<AcV7Zb_#.,WZ3Q9:6DV_8916MU=0
=1P&cBM6)B(FdO(Z6Tc:>)a?OZ)Z-X8;;S362K/ZB=c)4?EeM;Ga4g_@X<&g2&U:
@K^P7=S+FI9536ODG\f9UYLZS2]a)L94\S,GegK-1JF?&4JRf2(dfJ2=]2Z)HEO-
7<6_]cgF0\\QN4MdB6FM1?d#]A)YE1^,?WOFDb<CUgJ#dYW=/&>d(.8Yg46dZL\H
+?8-21F17>55:F?0cgJ6[3L[65FcNSP1(V25##;L6.^W5.#c=K),KZ@.f1G>1dgP
dO3I;d@KDN41>LZ+\La8ce5NLYESWb\SWa3^@@g0^]DcfZ&]@b/;W@]4TJSFQc@[
:@aXV85HR&\REU=TX/X[B_QV-(G7FITC[RXJALM(VQg@=KXACe4Ef.1=Y&#U>Re8
,?VL@QLNTUGf]:0ea9cRLYF.6ZS9\gQ^+IM[;,:.E,5+,N<GC6Fb(V:Nde^Z[(^:
>cGNNMTb6G17ObE6R6LD.>fJ5;aTF9VF&T_B,)QT3-C49J@=6[)UB-]7U&Q?C<a^
f-5A2RaA&6ON#]&I^CFJRfE0WP=e]T7_+a6(2V<K(V(<[-OdEV@N9Z)XR44X;g(X
DVUeeA-CWPPG3ETZe^)_Y&\)V9cH,]C3)7&1&0PI,3Idd:0&9b-(?]gO?NQ^CKY6
/MeB(-#De8eB&0^;AD;]DM^b9McYS>ROGAZ>2_R]2E;II2T_D[(>KB8&Pb;&PGO:
B4M9F8fWM,C]fM&1C^6JH<0Jd(O0CN=&\Y4QAG#?(A/YWWg25GZ<E=?_;g_]2bP7
?COGC24CY=QD40?4[b;V/NegFXX,7N0XH6f:]\B.JU=7N&56g2=\d:&EG,3cMAXN
A+9NU[Z/8;F_0T16^7[NF]>N\\&\d1HagJ\Lf\)TW-+WbSDCBF\4gO:8#JfW,<GD
O4Zffc]a9XEH=g49bC1=AHBg+bXOIZGcf5b9T2Q)OI?QI2\8HG)[d-4BdOR-I+A6
)C+4[P:e8,O]?E]L\a89HRb1[QS&68<^b-^g=eZQ\9C/YRA&#=Nd?(]_0(HWg>??
./8.?;[4fB2a;-e>7&J^f2d=D?(8-?ZbET1,V24EgWW#LNDJP?&a/V9LI2T]\72/
Q\4&N=EF^2YI&)c<G0::fZKRFc8L(b2/>eV-6_cTP7dFF&2VJW5N/<80WC71D#9Z
&QXFUH?5E\G3@D)#fTK&fLXg^Qe=f?]X]YUa8-4:G+g+FaP6N1eS/6QRSORP-A:@
3==_AJ_GN/ZWe/<2^MVf>D_#Lac;@B=UN(X,T><V8;>#ZdSS/e7LOIG-+;aX_HF@
d0R8.1W_Db,1A2]JHJE,<XCFXU\6W)>-(#._LZ2N)B]c??<C^6aM2+T#G22fP\SE
G-[<A.-fF&fNbI,E9],#,HJZ9aH1:XYdAY2>?/QHbf5B.#<,9faAd7e[1CSZ,8#/
K]P?2NO013FQF@9]3DH0_H_;@#ZV7-1>>C@U?c3(@OA+&TO6[PGETa)W7C0Mgf9:
466/d3R>W+Y^6M6,QM58DIcDXU9.WF^D-6<W-@(9(.5IDYe[4(S?BV)Y>G1>FU?A
;S##SH_>TVSY7DTfA?@afAgP=CZF#:)We_8OZ,>Tg1a8?MPeRQ\EQ=a6MWg#R5]7
ETILPN>dH]BHOPS#L?IU>YROT>f=<R^?1FJRXOB&OD:T7YG4D^VZddJ>bK\;P)?W
I:]Dc/K);SgQGXX?D=_<A9OILD;V+X4T;W];1aeQF3;D/^9JQW5=b&6aX5S76YZZ
/N@?Z1Ig<WXQXUIQ-.3I^>BWb[_5a79OHP&3Y#AB+,5B7fJ[G1SH=HO+<WUdG\-H
:/EKE,B;1K?V9P;&SEfaUO;4_)LfFP&2<NC+@_e&@YP@,8V/,?aU_?)D?39<]JP=
CW/562BGW^X83Wad2_]aFA_6KOce0MF(:6)/D?8>g-9Y3DQ#dS]II>59X,,7>+:R
5)]>E?;&#]beeeI(ad3f:c>2]HZV#(GPG4-]=e12ef.@T8>4;^cH?T(Ib4bGXT,(
[2NYP@Qb&abCAHIVG[1>-,/QI^#3]BXO[2V^e90#(^OBBL13DVeaCg+L#;-cGg.g
:W#TC2fgaFKR8g<KdLHDYd=MVPU>6).d5a]F4JPHbE^=4\-+2E@9F9EOd(VECON-
P6AUSE6TKPR3E>,W(A[/^\HZ.?\9:UbA-VMX#Mg6bPKYOKF^D7V32OL,9R5JR3Q)
F(CKT8[_Z(gT<-K:Te7K&e\/FeR94=(Q=?=Va3Fa?A70-,G7Of500N+(a<<8]L-?
@^U(KC^BR,>?fQ)HB2X8E-TbD(E\TP34F,MZd5+(S526ZZfWX^)(G,-@f+,?0?V<
2=:WO;II\e,4)5-U>K+dQ/Y:(C7TB^MfWa>3,]a?Z.M-ScYcH3Ib4)\5R0H31>Gd
VQTOTQ7NHT_QNGe5F3#d,CW^(9(P03EQ3MZ@5Ma<KQ6D,PH-DX,2gM=+;MMHR<_4
=+e23/A(R5a10bc>Ze:UZCU1_4&TR-@I^@@8+e#YEBE2TLJ3#a]XDB\HLSS)DET?
G(\bC=P,6NRS8dY3G;><D..9HC43::^SEDI=B((XDMc9@4[[@:WG1N?ZbgH-\6>D
3W:dAI+ZAbU9B_e^_-eFM>PVf1&_aNFH),V5P=@aXWJdN;>X[eIN+TAM#[4CgTW<
RH_DWc,@cOfWb737A@Q3a?0@XW^MI&aJVaQ.D]^93B\I=@-g]8UfW8Wgf-<&aT.e
d#^<8?1,6a7UH=8GcX<E1GP:T--A.a&K2/B6&\PTLVgSdOVf>O6Q5<2UaaW5#GFF
dZ,MP3Q>ObH2e4[SGRPGcc+457MVEO3^MWY;:]b+d+c7S5&Y^YSJ+5CUN:9,(H45
>4<FQ?(5B=acFC,fQ<__:B<WKaY4_Y8GQcM8-E@.3d3gZC^+W1>.c[GEB)+D?K:L
XPAU.Cd&GME354_dcdQ0Ee^<@B[S0BT8HaQM]9Y90PXV?K5J.dWO;^Z-63DLG[1F
dK+1H-;4Z>8W\-LNGa2Y)S:fY=.I<R2#Ta=[O)9b9>aRENKbG>0eBS-?b-B\:(Od
JH)_YX^deRZ=AB-I.X>VM8YN7?7EA3?O&/>]_O\a8c1EF5d17H])2G<H&T-BfT/_
T@I4:NIPR9,/VUO46f=974F(bX2I>#P@.)bb2HfK:[(TB4WIME-VB@2>O,MOVaI[
ICM5+e#Dc&(M?(>BPJ3&d9&FggW7[IR(C6AQYW4>LU;AHf5=V]X7=2]N?@,V(5],
3M4@PReA?VIOMd)dK1G98QFEgHJ.Eb[&>Ef4ON./-?J,TXH]7e\g_]ID,ZLZ[RC/
4V,f\C07U6DRKE&G@N;LDb2^V2WNUK100P8_Y1Gc<R5<[cIAS43U(&#^eBJRH6+(
SMNA\eJR.GGRF#=b=5/d4HECfJ1/cCGG<g1A^>>]1H]b/.KHFJ-HFfK&Hb]?J)MH
EHK+L@[6Td>O+WJT)+e3?C]M?C+<4f_=HI?D3,+9NUDI#Y\1DTP2VK2,\8cT\/7D
QZTCXQef,#MHc3FV19&-)H3ZQ6R:5@=T;=:F8/#NB6XOOV6V_5d[IJM[M><Ma#;T
@[CFE^=1Z:/H3@C=2)F:?1SJJVXJRCCIMN7,OdcIb^7<2UEQ4LN@J]HeO)K9OXVd
JL7cGa7I3>A8,+<O#)JOQ,@,GY6)OfX/E10FG4/A)@EfMNMT=RV:A:XT67W__TIM
UF>S^^?@&&e/#gGcZ(26JB4/41;D&(PEJ1G;Q87R;Wb_)P7:S2dc2O:0;B=WXWP1
fFSb4\efSZH_&NIC0[A-2=5E4SHVT9@.Y=]baZ-Q_f.-.-7WWUTOM-O89a=b8/+J
]^0^3N\#V0-<(ER+/1@XJQ7Y@Da?HOYDUbW7db-gW=dWU4M)fXgESae9B\&623#8
\f2ZVR:D+eP&:f,/<S>L#3UX0/J@)WWF#Q;YT77\,.E5)^e-M)PJ#XcSGP>(W-gS
A1^@]6<3/\,C4Q]./4K#)):J8&&,e#[Ba;:Sc+,>^23/9bE0-YJ,JGQ#W#,COU9)
YdJ5V)E@B8MT,>^L#ML=WRN_)3dO8)E;BU#IV:\a7@4c:bFKOaYSCU8_6WUW2O.=
NX3TXJC#3FNN+8^cYXc8<f>J@L^Oa0]6^g3-94ZK:)8ZRbJ64G\D\AQODXW1-gG^
S^L\-EI3@:STYPI\gD)7)-/?.UK+-XA9\;]b_&JfP+Q,YMf>&7>AZ7&UL]I[Q;(_
bef9@=\15D=cY6G,]8dYGO9XN@NM57Ec=JYZ\=ZC<\7Qd]DQJ)ebdVL6CedT(Tc_
6SbJ>JCaGU>U);X;V#DQ?-5aI-aBKD9:0+^5H]6XP+7UT<f(?),[9O)=(DHf6A3Q
W4VH:TVc\V(Z8/1ecG4(3BN#]A4M-0W\UH3DABSFdC&A,dVdUSVcC>MBL9Y2+C[^
db@>2>UYHIRZP>3TJD[_Za[dI)JBY?c5U1Z)F<8F[7R8X\ZNNg)X_HaERa4:^4-N
(R]2O6fbVUY#&A#@cTXK_;P:7+1<K5^)RC_-_fQM_=[BF##eYAPQX;dE0NJ[dJ)P
&/WGIO]1g-#PPObSY2QWSK4.H9J3&gZ7G@Y\aO,aES>AOIW)/3CIe/:IG+^I:fY7
;Z:3T>05_WQG>&PaYFd#9BT3\fNQ/#3ON?S\I3?RcZ:G(eS0E?=RV>8,AH-?ODBI
Xa4;:Q+QWA#0A)VZ,?U2b3S\PEJ-UY+IJ:]aWIZ?SdFIMB8DeP8^01]geC>&_c-a
B7Z&^>^>HPBF>?4WQF?GVJ.ZV-&,S&&,07C1]K7=_7NQ/4F8b]e2Md4(YTIQ9FS4
K=,&5Z4&aa3+[?OLA8;_b>8)U9IX,;539a6Y[N-CeB/47[1&E@J]cD:5@IM--1Q&
N6-I#g@55HETNYQO\8U3:&GN(L[H9:OTREORI#-H+20HQ^JY30B<AY1B8#=O3BLU
Bb]18Z(=2Q\ef6fa2d^gccb^O=?G/=,\>e^RdT+aa9+UIAVO==EZgdQ0,bN]?Y:F
_&\(G@/--A5AFL(G.L(;NR&B=YfEJfG=LMR5@aJ8]5\W+5C;TKC5KQC1,F]EdcJ8
XRA3])DCQZWF.4U>EH/)<FV09Q[;F#_>>//>N7/)YY24g(BbWH@\<\DO4f]Gb;4D
9EEUO)LT<0T#-(PXL@aZRQP-(#&IVR3IZ_V0-aK,O^-eY:f3fa==_Jg0Og(K/WM=
X5__&UJR^7c35>W/<WZ3L2f+a\7Z_?/ZNIW;c,ILO^7,WcK,.VAI0gIK/B;dJDO?
SFPdI>E1N)TG#);,Fe3:SG.?K,#.0#55[OS&T#bQ.YJPAL\4dGJ-H0U6O.QTNO4D
0J\TM[F\ded;Zf;;()fT@;,ZUU:aL1YI(21Dc2_U+\2D69\XV-:0<K?.[MYP1K[9
67fDf_B1W.FGJC[94gY6@B1[N@/-d^c:58]-EMCZ,9>5^35f=8S1ZfN,(DZA0c<4
Z>dUA7TC2X+9?Fb;RE7)P<f6=d]a71\g-K?Ne2]_H>(OL]CRLEee02gGC-(8g6Q+
A>0gf5R3DC,03UEB]U<5a26;9aLb6M3.c,9Y=O:X\XW<EU&.VA#KPVB#B.,[>Ide
;+KSVJKJT_TKWa^?IO;g4b\M>f7.(BRB5G[,=TQNI\BB\bX/VW6b<UeS/9gB7g4U
]T7@Nc#R#9_Q:e11V5?MVG9DU0^#0UJW)RBZ91-]fc[SMEf4Vg:B9(O);6K1LDW&
T;Mcg8@AM/#XH4(59T&GI:9<5C]=V=>KHc4\:f(YEF9XI2)6;&H7G)V#f?O;?Z\3
SE2_M08/ILM;d>.8QURB9_5P9Ga:<IY^;<a(LfD0:CeUUA574ORJNP))cS9=U>DM
S_DO^NZK>K?&?3KZPE+a,Dg568BB].g<dc\I0QQ3K5f8a7Q()=R;b,N,,K]c^D<-
VKB:gU]SdA?U=@1La)9J.HP21_0EVXZ0=P^8e\36(DY(Da1N-U2WO9)V9ATFGe3Q
FHZdQb>3X0[HPPPcJ+>]&W(Z>_c)L&gebPSIKSCf67dOBZ?dZ4,/J4(42\RKe>;@
37DWZ2P>8e_6CbP&eUR/#.X:DAQ97\&O>&50K#8[463Q^GWA4@#=#6>51Je[\+.Z
#bFGCg>;UVU0g@/OI8W:,_-^S<gZ6Q+Q+F&KdX5-#e-CTaH)UbJ&?P_3Y2@eg@=R
I-UPZBT.9;Gc2XB:Ug/@V-(M)8)8H]e8g&QCCA;U2gSCX&NQAA/M/U]L6XM5#HXF
3O2?;IYe4.TNUS+3\M8T/AA)(2gUF^g#Zg)2EJN<IH?dPR>8eN\<P4C&D7-a.Eeg
/Nf:H1e2]KIdF[201\<ffUXIf.3ALCF9Q\-/f>_8LJ4adcV<LF2CF6R27F)LNVCP
cdNJ0AV&LNeNV+IJLD9D8[c.MG&^f,.IMA+5?F&[_)SY/=U&TWC@&;-c()\@N[c)
6)\Y63A.-dGSTU<KdZ78M+YfQ)&__53F7UT#[#TZ=&cUM(FM,<:;5Jb]YC^88^N3
T3_.:<KL4T426G:.#Qf\e(f.]UTS#EF_<>bMFF@SXD\2J^T5P6O^;[V(&G=-#CQY
cP+;da&f\W-0dc@?D;YRWL8]NQB\]c[)5C=4V1gRTIHdG/Mc#T\OQYa>-S#Q0S/-
65f.,VIG2G[:a#Z&G-aTM\?JQ/bc\HJb)_<LMI0N5UYY)(;XI:J6M/dW3AX5_BYd
.eM+BJ:e@L1>^fL&6;Z5f=>9<?91>5;,;gKf,V2#4Qa4W-/cJceV/AEdgT5]G&@2
&B9[(7<458@P8_4&-(YgMUdQ1/D+U9K/[.0,O7O-6U6-MVSQIN6H[U+L3XZGG1Y1
@dV5aP:^;cfZU#2GWIfCDC>.@E6/2>9fLLY,Z,)K6(cbKbcMG#8_:-b?A?]R@EPN
]?E9#G<#f++f[gD+R=XKfX?3^+[YT]f:EM\,J#Y\N[E?ga]4ZI>M=(3W?C<-6_EQ
5[-.;f/2Rd#d7UUKO9K,Q1b315PUQZ1A;UPN36E9J=)KU,5@;<>BD)^Q#>5IO;(2
W?E:M<Y:^MYH)I;Bc736B#IbB41OTW]<HP0L@L;(D\E[;-N_Xe,6:Z#7gLZ02Vf4
6M:,C9@YJI./)WYc/Z4)6M8/&d,d70e5864<IZfD/TC1bR.bP<]<6H>IGY4U[F:Y
-P:.,^+WRgCRW<KQEQf<[8JfUBf6aM?JcNNd?c?Q0+cO)676V(4?TaIc6gE;?U^Y
8[F+[7_G;GeMC8WIgMFRR\(.NWXe(_4U(/9CC,Vfd0-FNEMLDNYd.#3EO>I?0KeY
^TF(G=Z^>(Y,/_.d.4]G7_2Y22GL:>QG2N8e0A[4;8]>(+3[D^I+UU.#48Mg-1UY
K[d\E/Z.(32]LE,W.:THd_HgIU]19N8VD6LP7V9EFb6[R1ae2BAUHXWJf/_AUdc-
b&](,Y=bPIf\;EH0BW/Ie=/[J.,DR9SY[5eO8=,Ze+aL-bPR24bZS8#F/S+OAG<>
,\A=(3@..67V<fg5-.0/QGDBVH^9_6-KJO>[2^6X.>OVTF_K>7)S\gL4PHSe=;QW
Ve4?#WO_Te+9OFX?>(EEc<TL:F(IZ;T]63TM0gK_8:3;_dEQ8Qa3WaEA^69(32,\
g[<dLN2QVcR\&Db3b59PG;cLJ9:abLWJ9g0N6;FXF>Hf]e1:+e.DCKb0GYYX<Ef+
@F^I:K^&8A5-L+S]#J_OY\1,A66,MTc5HMb,4CF(-+OWg66c?S>=JO_CKB)a38F(
C,X?BMU27^VI2LS,_EL6W_4YOJ<)SWI74TZe^f#1@[GS>(3Q].E8<6DL\JL450:V
:)@->-G7M<dX5Z#:84DDcBD_3R5+,ZTLY\1L_=A^S?F,&PY,Hg+[SO:#eSQb[+@R
Bb^O1R.b,@-,:dU6TZe8>2[cf/&4GU1e4_W6c(-J_1dEIA9&X@(2,bA-/(aQY/aB
7?(^O9Q8dc7M^;LT>b//BI:XfGG+N=&XX>+E<L5<UB34X2+\CV5#3eL.1(U:\8aN
VXd.@#cB_.Fe?_;W9BT#8ad72EeZI4FO0T6^gQ\_S3-3F8/7_)<KeSAX-<bJA9^K
\CT.69SJQ^E4:+I&EBJM6b:>UP5gDR]H]1S:We36TNT]L@#/>,B7C^PWcfA:NXf-
L8b7\ITEN^I;aCX@3NFbFJW-WO^3S8KaR99eTQ8Cc]78d[Ab^?I\D:03X&c3Z+4H
2]M8@/_W-+]R(1g5+3gD\,,SgO(9,:TcJg#8C=,/W7#]MOb@A>\)(d4,8#<&FPNc
eP[4&Z(DaLLE:#SL8f(,BT31OGF9f&<VE;-M+J9Y+b:aMZT4f>IDaH=.g-(1=dI?
CR3B.@OZ5GP-V,#T1FaJ.M4;4eTdRgc_M7Q.J._O[e.LJ>C&FOaAdNQ8^_R31g0Z
A-)1Y#2cZ2KCW@\DeD5+#JeJ0N,H8Q,/5TFVKMN,+(-LTGSIHa?cLUOJ/ZW2QbX7
96g-^.40_K\)-K[<TI\Y&FZEg-RfM],9MLeea18]c9Hb7M.2R?Oc0Vf2aJ:3agJI
.gJ@&EOGMOAY&ZADP\KB3:_?=@K+:#RHIW+/YR]gB?);.dQg:cg/N]&ZZ;K552WB
1Q&S=S)[(H,\f^9PL:;[8=?PNF1TJ3]GK>c=XgM=FJ\KfJJT4:RZXE>cL,22Q1_K
Y?f@D#\ZTZc2J<_,)1YZAQJQ3?]TFa9H(.aWZP[+I3)82MAb&[UA1KA0VeXV4Dg_
4J>&\B?1D[dfTZ,A0J/:&]DT+L2E^.#1(+TSI>1:8&#=gX8e7AC]2#-[T-cS-OQG
#KY&^AgdJ?:W(&I\+aFeP&;48JfcMaU6N@)aKX[DgZT[1E6UXJ)OKGE,25D+W2b9
+;d@;g#]+XP(R+3L?0AV+g4^:^>=Z+<cb#0ZD6LYWFc-0F<LQbM\R[(&H0;b/G,R
,O)7U=P_8\e^A,PMXNBB6e9a\DL(UUgc&[=g:M:DRQ]/ROF[0?\RVF.fa+#UMb,Y
:+S:\:^aK(.eS5.G,&g:[ZX>XbUN<Mg:^A&A:5ZH4RZcAOW0B59GP^2CMF.K?C&J
N34053S?^PX;XF(R-B?X&;B/^>Of7DUJ11?ZJU3MM&QL<BgXJ;f/?76_dROQ3[DP
&ETW:J\@^MU#7g@&4bZG?;A918OWQY8G_fZJ5(,[2.(-P().,c>TR-Wc,8#fDRIS
5dI3c7d(Z^Rf_NZI3UBM2JOXT#aBXKa\UNgJ_C=V=66BL4>0-J,cT.W:TP.ML^,8
1<X+3XF0IB2DE1]P4b=?Vb.K>=Xd6?]3^X1([+UG8^0\ee+?6A#HU5,/EBa7;3GE
3V::?g6Ra1/LBd,WCD@^Y-PJaA95+3H=^<S+c1.UXK9MAce&FZ<g?TGT6/TOQ#T\
JIT)XMF+:J\M87bJT/a_9c\<4(;Fb[ICW._/5>I7&4O=KREbG,TA4BHP/J)UH&VX
_/U3Sc-N0ZRVE]3^QW?WT?cb+I]D2A\WHEHF]Qc6F3b\H;O&0BC(3JL/D.cNL=X5
JK7M)E:5IgR8UNFg1@^(cR=WC>dNf\.C]gNKg&?&&9N5J&G4J+9Z,U^2/Z8^>5]+
DggPTZe@.5OdX7=;PaFM?_(PXFW93[>+&8WR.P0QXZ,K17BI+9aZRL[FCBTHZc53
Z4c9<;F[+\1F<MQ3CgN#>d>RO;bK&P6MQ\T)F\;UB#FeUB7)#[ATI[M:.505>[@)
e66W(=abKJC4Oca(:O\4b6APUI+V+_C?QfU9[Nc9#Ne#Z/Zc>/,ERLQ[6T3_,CAJ
aJYGd/U=eE_2fY4>7I?gd6(3NYc7CDORK>O]-[()=^L/FEXHZJVbM_>935UdH\9Z
L:JV9E+8Z6e+31T;C/e9?P4X[d1#MV>gT#DaQBg([Y?W^>YW,Fa\[HQ<XR1VdJ(,
QdR?X=41,.76]<(O.Ub[^T=BJO8=W[LB#\8QAB9V<JI@?+]F7<cY^b>7OYDX0b@X
PcJM:,Ue2gS4DEVPg<eY0IV,cOCM-e#VIZ8?9M6#>]NB\Df^@]4dZL<=F0JN2WJS
f]?WUERa[c77;O@QY@3OU-bbOT)7:[SGeW\B[3Wf+2<ag51K][25P0H,dH9)dAS:
U:-A#8,@86#QJ>LT=W]<,[DT&dQb?cI)L/LR-E]K]LA<W;54R\84@7<Y&QU@3f>5
=&S405g/.1NRA1.S&G[W_OV9Q?cV@4(Z/8Xd-RU<0Z/;W_c_c&N7e^-1+ZdJ367\
\1)Z#=\gF[YDQQK<,F;aRP^&cO^MCUB?>RR\2C,SQVL2UULAT83#>E46/&V&+NX@
3+Hf99\I)89Kg4]FRV8^<eL-d][g4eO3T_#Q)&E;\(P1RO8WW9B5QXI>b)F5DDUN
0H[0R>VU]>OLeEJ9D2BWgc>29g_=/[cUcX^.Od:<f0eA.9?3-fg)7:ZU9fC/YG(Y
;ONFKe<J1-ET8VQ;M9\RS)YM0H_.6=<Bc+=I@9LW+L6gDDT3QB9Q9G+?;P_@B\45
K^UedV1N=fb9&2c2653-EU_K0-6/D1LE\Z65H/aPF1H(7)AM&9AYNaFgXU<-_.#G
ZK[.AF1^EH#NL/U2+P#Ff?^[6IX;;,G\,KZY#g<,74?F<B>&0?a0[UUN7)afLXGE
9eQTPQR0G50@Y@8]_2g8EZI?/)O?KAY5S.V.99[M@_#H6>V4Wf-@<X\7aV<=STFT
ZeKfJ\fd>K5,?2JaND)&/[0-Z=d>:]cMVf5U:W0:UF)gQ14V/F_M.CZNCM=[d?=7
2OT4N4XN3Ycg2YPWJ-fK]6N#(+ZO/WFd^5+cLc2-F^D6aG\Xe<73P/<R1H/L:WDT
g1gEX+YQg06ACT)PHYY8PaJII++F&cO[L=TF5=\VP[5&E:;GJDP+K<NCBQ4\KX8K
^](f984M-0+JES>T;MHZE+U@eR^067Dg14;XCccI;2DIJa?D@9F5T-GRCbLYKT>C
];(g1LFF4LB2TZg<ZCHS;RPaU651a9D;JLDdg^40#2,>^>bM?I^#ICZ8C1CWf.U,
V+c.6<HD?QK3dge3DC7T+0c<->T5e1T,=#.dM0d?)VEJ-Q;#I7L3XZOFeGL)7ZYH
U-/F,2TR6S,P9A9HdQ7eg^P&K)d4KT.-&8WSSZJTWIb<;+H1Sf84B<]3U#.f>_&K
;2@3dMJR<eZ].Zd46=H5[YZW/3J7G@H(CBJ^\:ZYQb)1A[@L>O0H2_>=_@M<-LBT
MD6]?VWdf4FH8??Ef[V5PC9-&dYCL/1ee0dB=-(g>-_#<BGK?3_]HC8e@IH(1H1P
X^(XC<@S2U,dGNT7/(JK@1@bg4(:Za:Lb#gc5EWXM(&MWE#86@R<7K>cMFIeRC5.
(QU\]AR-_.e;TBJ1+6R])F2]??[OQ]NU7-@>ZTALc[2#NL)[))?K6B@Y+=Qg_-ED
Rd(H(9fF\/\<R]e>,2-HXJ0FT>.3/?,:V2BJ(OA/K_CB1N-5TC\T]0@6.[\,6/Gf
D8IV>=[(HZD.g-GK\fEDL[;NBGeFX1DF4(H62R;3eAK(6D:NUPf>XE#(@0?BTY+X
7=E=&OKR(X<Q+[Y)T_ILK,ba1F6TGZG@FU/>.c02[-2S\f,B\eX:9-WGBBYR2:)_
-L8+gSH-/3A:B.OOI[L.@X1GM)L=F&5gQ(?E8aA2YDHaGU\B29H=LB0JbB+.&]_6
NAK&[eI[,K7OAE]YF>5<RVUWH_<,38#NW;O=c^6)FS(@2c-,)M93#(8bRbM8A]\\
L:Z_a0VKJa->OFc6IG,fad;3BA_S767J^1/Qf]C8ZZfI,>gXC9E+[GN:\e.1UcIN
Nd?4e-62(,_B5TNU;^+MHRLMLA[[XYe_DE3]J(MLK)>)VR06JX:#+b3FcX^+c.3.
++HC#Lc)g&.9f&M#Z2ZD.:cY_7&=P.Ebe4fD+,XJ4=fcd&3d^Y0[<8209DH^J62\
RJe1b>9GJJ[g67RC.HRH&0_efZ#//Hef(a#a+#,d1H_SN7D]^0-)UGWUCFAQJHQF
.?>O:OVNO7ag18L\aSE_9Q)N/G@c)+;(G:eV.@O8+ZDb]U)_(_d9DZL2FW8N#d[@
TZeb4ZK/HKAf(QJ+PSZ\[#6Ga2gWaDfN.@NPE57IP/&eQg:#,[Vf;9aD^)4e3<a3
dM7O:1N)[+N]cF9STaCM-Ya0L@\=Y<XR58AEed:WEVZDZL9@:JQPHKWJFeaL=V,C
Y=Ff;--f[Le,7gFJ[AY1C;(FE4]Q&TT(M9,0Tb)Q@BZYDPa8#bdY3W_^I0[ZH3FE
Z?CE9^TRM_L+B8ead]#?AQ:QXW]RWM[I5FecaTB\UcZFaIKcZ<V+VD?Y]AYN\@;1
_.<NC3Ic1g#FRRN,.b:?:SP-7TUW/db0\e.,60K]F;8-06eI?g5HMe&6.Gf5:<E^
W9[Ecb/Hc@WW#WEB4IVWJMe47,5L_;D22Z/Q<2=B^g_EcE<;S4;7dUeYHgG_c9B<
4)&.gTf@=2c[D.@4_.-BK9\FUT\ZP1>C(1_E0]fB)IRB\:HS,DUHM.FBT31W9/PT
D\@.PE7L_@.BbK8U:O#gFfEXE\[I#1AZ9/++NEJeK47F2[C?EON1S=4#KeF@@K):
g7(2,c4Z>\(?g(\1Z@?[?b[85aPMR8I0L#e5_M[Q\M,P2U)74cN#KdSWDY?e+X>S
T/N9&O3fRUY=f.6XB.NAOMI)(M2F]KWY@b:gK&J0gD+-(Iac.Dgd8V1WP=I3>=2V
)#1</Z.2,139HG@VcZ>A1&A(Qe3F=CgQ\c@dOD>(9W+/^L3A/<@10VL=M>&9<(4b
BD?[X-f+(L(U=)=;ge1RO7<EMH;3R4A#QZa?]@^D2><46]:g_6^.4NJfFBN<T5@c
W\1<.dYL[4MA&,:NS2NMB,>;RS9Y[BG2?<PcU4?b.6;,7gZ9TVU&-\gF+-X?_.17
14#P8Wc99H&b?=P=QC4)dLVM9_E(L[3(B]J(),B-6A3?5e.+M3;#d]AT\&bFaM4B
Y65V.)C9^(DH>.GK]X=)BSA5cH^WPL5JP)#>364TNHeG-O]>?e>7=9X@U#XJD;[F
?PfWRbHT43]?(gOM8(E1d^>G^f\;DT6DE6MN_^>=K&.[[6Cg1B4;MC>++JVTaR#Y
C7QE2aI3M8I3:R,ffOTWgUJ@;<1/bA@&.)6ff5;\_O/K40#C\)TU]XLG99#9c1>#
[&,HJQJJf?cg?M9^fTC,bVR7_Z+7ISRN:a-SO3LK?C]7b)N/gR-QZd,gPY]L>4dV
_e88;8Q+e4+_2H(LW&C2PU..?=S-Z2+/CEYZ]T?;VTaS656D[=7eQDb_)?5-e8V(
MFD3;Xc4+Q/X16U,ed5;R\)0,2K[QOP,@A^E3b>G\dK3MTODb<3_)D<@3ef?&/AD
UI1Lb@FZ76HV4<0E-+<g2MJ->7SO9Y)E@9)G?IG43/#6);_@f+,<(O[BY3d_XT[9
b^)cR.(DL4PJH\EO0JA3QF:Jd<O.Ge&cb+2Y^));VWZ=)X/&H0A;/.bI)(M95:R]
=8IZdN@KTcAOVA:fS4ZcK9ba15H&Q+FI)(M3\,>1gJYe]]6ZJQ8]gaY,O0[()50d
fK(E\B]64I<X[2)3V8D^&1R+K7[D2QbMU&7-^_[f)e37&,>^>-)/_C26bA)L?EE\
]D]Y=FOG<H?LcaKC-]NP)La+;^:)\>=<=L]OJ&(;IAI+d]&cJ]bN<A9O1?;\e8(5
P)3HCIC.DIJ:fIcFLAcT&)<Q#2&c+<g(IR0b(VOa\L+FFFY)H;J>4,#;-C7/[fQb
5eV=M4033Jc62D)CfHVG6N,QeeL[S58-?6FWPIG6.;1c8RI1O((@[.;691g?YXO7
Uc3NM=&-Q?4PQQ<T?@QD=LXTfge4L1G8^7.5Y&Ae1&.71&WeWYV@924f;d;P??)(
(EEV.3BR5KO/)X#P1eI;>K<3]=T5<^C?>]/C0AJRUa)#c##SXaW))<DDFIB-OE-L
JFD:CC@T?\2ReKQgDX@MG+g?a(\:DN>B2@XdZ;/bK8_)d;UD<//?9=BABWdSPZGa
2d--fGb3@]=PT]=<(:9^[OYG6.e^K?fQF#N9UMAU^2TMBO3.D7YT#L=1+C/E&56.
FW;eGgEQSfEPZd,=RcDBc7\c@WYX,+?<BQ&;Xef3QDE3gf0fWJ.G;bW+N_e=N<]O
;cc]^/]QJVdYB5Y#7\?YL)]);R-A?UNF#)W1;2RSP8@_f^->)BZ[&;Ec1<<3c7)R
=fc@@VQ+bfW]@/RDX_93ES7:TNcT5S^ag@-LKZdQ5>>/1)d/bS.bBF\AGCIGD;MQ
,5+NP)\WU#I(WVU:,T[<:?GBP&]23NWDOVXafNU040[H-[3N.(RD[,X3DUWG?/Ug
5EfOPdcO6b)^4;be\&FZ:&g4Q3N?:>?X)3a?UEPA2=T5VEC?4f8EMEV]Q5><7W_]
R,U].6gdbD5HWO2cg4Q?9d(MH)MTPA>.3\YfS7L9bNXR9^SM52)gCC8d,@8IR>N^
b97)aQN]R(F.VcQa_gU#AG4#+cb_)E9LSJNO69fUdZ)[91S?_72^YQVY#/5SUXFV
WZ?[JGJXcB/GDO@gbbIf<6]W/C_-]HS)LLaF?:[VaK23(&/T6?TaX[Dad0PQON5T
D2II@K)48OZ]MG8096V7JGV^,)bOG;3/d(B][U,[)BB2>d?M>Z^8]d(b5?AA[Cce
L(<I&0^&#c^\=\#f_AB&5b-KH)RO]bRAP<M4#0&dO5,LTAaLE>HTV8Xfebf/W#dY
@YL#R+/B_/Y8KJ)-17VcPBTG\DL4]U^UUCb/dR(377:KZN@K,.:EKAR;@/X&H>&V
dTM;1V6acU-^XQ@=T]0<XT/B+-a63.#9_RB:&BP+4C5OF66L8OeCYRN7N#V9I\RE
9JB#^9](:><UYHX3B21)fc5UYUSF\b)?L=I0V#:Ee_D\2G+Q1c-,eSffc>gHe(3V
/^9TH7N?@R6]54CQ.aLV.]JBL67X-Dd07E:RZK8^0/F=T#_OUM1-ETK8MEKTQRe]
Mg8/OebJT;#Nd\-0#6Z\1#(N5I1S^RF_H;P-XC3]8G@YEJEc&<W/OT2@-dH<N[f9
BdAXW61\BKZT=,6@/@ST,XRHR#,4eMHaT.][de)cN8A203OL04JFR>+&XY(1KZbK
+>>BIG7ARJ6H_f\MK+@=cH5@;/7(&E2>>;MMMBWQ64F331#WQAS#MfeZd-Qa?5S2
VUSNO\d?^=7FX,LQ,>Q,a>[_I3&cdMT4\#A-^Z:\V-13_/OWS>E=>eFSK=K;DOW^
/-V]R_AMb7C>CS2W25ZSc-(.a\bdaKS;?#B4b8SP]K=47S[+HUT]KG^(Z3K8(T1@
DAUA?A<3IdRD;Pd#,;</NS/Jc\3APFUS7\6\C..^4W@46]LE)[JMN/Ed:Q(Nd#>?
0X6N]=gaJ2D.T/#?S_3V9CI+,W:gW#24&+cH8RN.f(f&;J\PNc,-\56CPb_LD-=9
)I^5BJ8+5Y[>gcBGEHWb##RMEgY,W[/d50I7&X=;PM_P.eba\Ac=XJ]5@58+T/eE
62\NJ:4;LbC6X\c9geBAW]VaE=GC]3C>6I#BD[S0TR?X;J0K+,^85:D\J\Hb8BQD
VaH;2CfeaT=M7PS\LF<g9KME;@Y^:]Nd(H=:L)RR7:\EWDDHHZ:L-UJE48f#;T)d
X9b:(DQ#DcBU/HDeDbBORP+GCZ^GIA4JRW7K,MdSUA-aXHF-dJb7M7(.Cab2&_f.
708;cL1]&-:3G??@2OcN8KW=aG0b[C-83&d3ag@]cAfJ:ML\CN52c>8f-/Y&NALM
PQ/ZKa)a[cM4YF<F:^+4@Ff&(5DU->[K;9,dbH\X1<<3KYEedV_/f1?[?/TIQY=0
A=?\4T6X3EVDI6)J(9F@<XeYH5:ESI[T4WeJ,+#VD7(]5+S.g385=(@=9&Tf?VAb
b<4&<U@4c38207F;gO0TIW[JgW&-_QN9OG[5(&g[A0E8<0F?I5aMXcAbU\AMMg?N
2O<7J/:M<_2XWBK6H-;#2B52[1GDf[&B:,QD2_W#U1Q>ZHJY>aS[^^,&KHY(9KI3
>g^:37S(b-bdL+O:_bON,f2Kg]PbBL-/GDUb3O=AdKX?YQ&C1U\\\bf97G;-0&E:
7@L&X/GR30K[e5g6KKM@KO554I-,.;\,9^b7[]6/?/B(KFbN,cNbV[P]g1GU(;BL
Kef+IH/Y9#T>WB=:FN5W\3:fd8N22cce]>[<>^&Z+1QJ.M&XUQ7]&6URL+V^(]e>W$
`endprotected
endmodule